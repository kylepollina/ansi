// colo256.v

module colo

pub fn rgb(r int, g int, b int, input string) string {
	return "\x1b[38;2;${r};${g};${b}m${input}\x1b[0m"
}

pub fn on_rgb(r int, g int, b int, input string) string {
	return "\x1b[48;2;${r};${g};${b}m${input}\x1b[0m"
}

// 256 bit foreground colour
pub fn red2(input string) string { return "\x1b[38;2;237;0;0m${input}\x1b[0m" }
pub fn red3(input string) string { return "\x1b[38;2;204;0;0m${input}\x1b[0m" }
pub fn snow(input string) string { return "\x1b[38;2;255;249;249m${input}\x1b[0m" }
pub fn snow2(input string) string { return "\x1b[38;2;237;232;232m${input}\x1b[0m" }
pub fn snow3(input string) string { return "\x1b[38;2;204;198;198m${input}\x1b[0m" }
pub fn snow4(input string) string { return "\x1b[38;2;137;135;135m${input}\x1b[0m" }
pub fn brown(input string) string { return "\x1b[38;2;163;40;40m${input}\x1b[0m" }
pub fn brown1(input string) string { return "\x1b[38;2;255;63;63m${input}\x1b[0m" }
pub fn brown2(input string) string { return "\x1b[38;2;237;58;58m${input}\x1b[0m" }
pub fn brown3(input string) string { return "\x1b[38;2;204;51;51m${input}\x1b[0m" }
pub fn brown4(input string) string { return "\x1b[38;2;137;33;33m${input}\x1b[0m" }
pub fn darkred(input string) string { return "\x1b[38;2;137;0;0m${input}\x1b[0m" }
pub fn indianred(input string) string { return "\x1b[38;2;204;91;91m${input}\x1b[0m" }
pub fn indianred1(input string) string { return "\x1b[38;2;255;104;104m${input}\x1b[0m" }
pub fn indianred2(input string) string { return "\x1b[38;2;237;96;96m${input}\x1b[0m" }
pub fn indianred3(input string) string { return "\x1b[38;2;204;84;84m${input}\x1b[0m" }
pub fn indianred4(input string) string { return "\x1b[38;2;137;56;56m${input}\x1b[0m" }
pub fn firebrick(input string) string { return "\x1b[38;2;175;33;33m${input}\x1b[0m" }
pub fn firebrick1(input string) string { return "\x1b[38;2;255;45;45m${input}\x1b[0m" }
pub fn firebrick2(input string) string { return "\x1b[38;2;237;43;43m${input}\x1b[0m" }
pub fn firebrick3(input string) string { return "\x1b[38;2;204;35;35m${input}\x1b[0m" }
pub fn firebrick4(input string) string { return "\x1b[38;2;137;25;25m${input}\x1b[0m" }
pub fn webmaroon(input string) string { return "\x1b[38;2;127;0;0m${input}\x1b[0m" }
pub fn rosybrown(input string) string { return "\x1b[38;2;186;142;142m${input}\x1b[0m" }
pub fn rosybrown1(input string) string { return "\x1b[38;2;255;191;191m${input}\x1b[0m" }
pub fn rosybrown2(input string) string { return "\x1b[38;2;237;178;178m${input}\x1b[0m" }
pub fn rosybrown3(input string) string { return "\x1b[38;2;204;153;153m${input}\x1b[0m" }
pub fn rosybrown4(input string) string { return "\x1b[38;2;137;104;104m${input}\x1b[0m" }
pub fn lightcoral(input string) string { return "\x1b[38;2;239;127;127m${input}\x1b[0m" }
pub fn salmon(input string) string { return "\x1b[38;2;249;127;112m${input}\x1b[0m" }
pub fn mistyrose(input string) string { return "\x1b[38;2;255;226;224m${input}\x1b[0m" }
pub fn mistyrose2(input string) string { return "\x1b[38;2;237;211;209m${input}\x1b[0m" }
pub fn mistyrose3(input string) string { return "\x1b[38;2;204;181;181m${input}\x1b[0m" }
pub fn coral1(input string) string { return "\x1b[38;2;255;112;84m${input}\x1b[0m" }
pub fn coral2(input string) string { return "\x1b[38;2;237;104;79m${input}\x1b[0m" }
pub fn coral3(input string) string { return "\x1b[38;2;204;89;68m${input}\x1b[0m" }
pub fn coral4(input string) string { return "\x1b[38;2;137;61;45m${input}\x1b[0m" }
pub fn tomato(input string) string { return "\x1b[38;2;255;96;68m${input}\x1b[0m" }
pub fn tomato2(input string) string { return "\x1b[38;2;237;91;63m${input}\x1b[0m" }
pub fn tomato3(input string) string { return "\x1b[38;2;204;79;56m${input}\x1b[0m" }
pub fn tomato4(input string) string { return "\x1b[38;2;137;53;35m${input}\x1b[0m" }
pub fn mistyrose4(input string) string { return "\x1b[38;2;137;124;122m${input}\x1b[0m" }
pub fn salmon1(input string) string { return "\x1b[38;2;255;137;104m${input}\x1b[0m" }
pub fn salmon2(input string) string { return "\x1b[38;2;237;130;96m${input}\x1b[0m" }
pub fn salmon3(input string) string { return "\x1b[38;2;204;109;81m${input}\x1b[0m" }
pub fn salmon4(input string) string { return "\x1b[38;2;137;73;56m${input}\x1b[0m" }
pub fn coral(input string) string { return "\x1b[38;2;255;124;79m${input}\x1b[0m" }
pub fn orangered(input string) string { return "\x1b[38;2;255;68;0m${input}\x1b[0m" }
pub fn orangered2(input string) string { return "\x1b[38;2;237;63;0m${input}\x1b[0m" }
pub fn orangered3(input string) string { return "\x1b[38;2;204;53;0m${input}\x1b[0m" }
pub fn orangered4(input string) string { return "\x1b[38;2;137;35;0m${input}\x1b[0m" }
pub fn darksalmon(input string) string { return "\x1b[38;2;232;147;119m${input}\x1b[0m" }
pub fn lightsalmon(input string) string { return "\x1b[38;2;255;158;119m${input}\x1b[0m" }
pub fn lightsalmon2(input string) string { return "\x1b[38;2;237;147;112m${input}\x1b[0m" }
pub fn lightsalmon3(input string) string { return "\x1b[38;2;204;127;96m${input}\x1b[0m" }
pub fn lightsalmon4(input string) string { return "\x1b[38;2;137;86;63m${input}\x1b[0m" }
pub fn sienna(input string) string { return "\x1b[38;2;158;81;43m${input}\x1b[0m" }
pub fn sienna1(input string) string { return "\x1b[38;2;255;130;68m${input}\x1b[0m" }
pub fn sienna2(input string) string { return "\x1b[38;2;237;119;63m${input}\x1b[0m" }
pub fn sienna3(input string) string { return "\x1b[38;2;204;102;56m${input}\x1b[0m" }
pub fn sienna4(input string) string { return "\x1b[38;2;137;68;35m${input}\x1b[0m" }
pub fn seashell(input string) string { return "\x1b[38;2;255;244;237m${input}\x1b[0m" }
pub fn chocolate(input string) string { return "\x1b[38;2;209;104;28m${input}\x1b[0m" }
pub fn chocolate1(input string) string { return "\x1b[38;2;255;124;35m${input}\x1b[0m" }
pub fn chocolate2(input string) string { return "\x1b[38;2;237;117;30m${input}\x1b[0m" }
pub fn chocolate3(input string) string { return "\x1b[38;2;204;102;28m${input}\x1b[0m" }
pub fn chocolate4(input string) string { return "\x1b[38;2;137;68;17m${input}\x1b[0m" }
pub fn seashell2(input string) string { return "\x1b[38;2;237;226;221m${input}\x1b[0m" }
pub fn seashell3(input string) string { return "\x1b[38;2;204;196;188m${input}\x1b[0m" }
pub fn seashell4(input string) string { return "\x1b[38;2;137;132;130m${input}\x1b[0m" }
pub fn peachpuff(input string) string { return "\x1b[38;2;255;216;183m${input}\x1b[0m" }
pub fn peachpuff2(input string) string { return "\x1b[38;2;237;201;170m${input}\x1b[0m" }
pub fn peachpuff3(input string) string { return "\x1b[38;2;204;173;147m${input}\x1b[0m" }
pub fn peachpuff4(input string) string { return "\x1b[38;2;137;117;99m${input}\x1b[0m" }
pub fn sandybrown(input string) string { return "\x1b[38;2;242;163;94m${input}\x1b[0m" }
pub fn tan1(input string) string { return "\x1b[38;2;255;163;79m${input}\x1b[0m" }
pub fn tan2(input string) string { return "\x1b[38;2;237;153;71m${input}\x1b[0m" }
pub fn tan4(input string) string { return "\x1b[38;2;137;89;40m${input}\x1b[0m" }
pub fn peru(input string) string { return "\x1b[38;2;204;132;61m${input}\x1b[0m" }
pub fn linen(input string) string { return "\x1b[38;2;249;239;229m${input}\x1b[0m" }
pub fn bisque3(input string) string { return "\x1b[38;2;204;181;158m${input}\x1b[0m" }
pub fn darkorange1(input string) string { return "\x1b[38;2;255;124;0m${input}\x1b[0m" }
pub fn darkorange2(input string) string { return "\x1b[38;2;237;117;0m${input}\x1b[0m" }
pub fn darkorange3(input string) string { return "\x1b[38;2;204;102;0m${input}\x1b[0m" }
pub fn darkorange4(input string) string { return "\x1b[38;2;137;68;0m${input}\x1b[0m" }
pub fn tan(input string) string { return "\x1b[38;2;209;178;137m${input}\x1b[0m" }
pub fn bisque(input string) string { return "\x1b[38;2;255;226;193m${input}\x1b[0m" }
pub fn bisque2(input string) string { return "\x1b[38;2;237;211;181m${input}\x1b[0m" }
pub fn bisque4(input string) string { return "\x1b[38;2;137;124;107m${input}\x1b[0m" }
pub fn burlywood(input string) string { return "\x1b[38;2;221;183;132m${input}\x1b[0m" }
pub fn burlywood1(input string) string { return "\x1b[38;2;255;209;153m${input}\x1b[0m" }
pub fn burlywood2(input string) string { return "\x1b[38;2;237;196;142m${input}\x1b[0m" }
pub fn burlywood3(input string) string { return "\x1b[38;2;204;168;124m${input}\x1b[0m" }
pub fn burlywood4(input string) string { return "\x1b[38;2;137;114;84m${input}\x1b[0m" }
pub fn darkorange(input string) string { return "\x1b[38;2;255;137;0m${input}\x1b[0m" }
pub fn navajowhite(input string) string { return "\x1b[38;2;255;221;170m${input}\x1b[0m" }
pub fn navajowhite2(input string) string { return "\x1b[38;2;237;206;160m${input}\x1b[0m" }
pub fn antiquewhite(input string) string { return "\x1b[38;2;249;234;214m${input}\x1b[0m" }
pub fn antiquewhite1(input string) string { return "\x1b[38;2;255;237;216m${input}\x1b[0m" }
pub fn antiquewhite2(input string) string { return "\x1b[38;2;237;221;204m${input}\x1b[0m" }
pub fn antiquewhite3(input string) string { return "\x1b[38;2;204;191;175m${input}\x1b[0m" }
pub fn antiquewhite4(input string) string { return "\x1b[38;2;137;130;119m${input}\x1b[0m" }
pub fn wheat(input string) string { return "\x1b[38;2;244;221;178m${input}\x1b[0m" }
pub fn wheat1(input string) string { return "\x1b[38;2;255;229;183m${input}\x1b[0m" }
pub fn wheat2(input string) string { return "\x1b[38;2;237;214;173m${input}\x1b[0m" }
pub fn wheat3(input string) string { return "\x1b[38;2;204;183;147m${input}\x1b[0m" }
pub fn wheat4(input string) string { return "\x1b[38;2;137;124;102m${input}\x1b[0m" }
pub fn orange(input string) string { return "\x1b[38;2;255;163;0m${input}\x1b[0m" }
pub fn orange2(input string) string { return "\x1b[38;2;237;153;0m${input}\x1b[0m" }
pub fn orange3(input string) string { return "\x1b[38;2;204;132;0m${input}\x1b[0m" }
pub fn orange4(input string) string { return "\x1b[38;2;137;89;0m${input}\x1b[0m" }
pub fn oldlace(input string) string { return "\x1b[38;2;252;244;229m${input}\x1b[0m" }
pub fn moccasin(input string) string { return "\x1b[38;2;255;226;181m${input}\x1b[0m" }
pub fn papayawhip(input string) string { return "\x1b[38;2;255;237;211m${input}\x1b[0m" }
pub fn navajowhite3(input string) string { return "\x1b[38;2;204;178;137m${input}\x1b[0m" }
pub fn navajowhite4(input string) string { return "\x1b[38;2;137;119;91m${input}\x1b[0m" }
pub fn blanchedalmond(input string) string { return "\x1b[38;2;255;234;204m${input}\x1b[0m" }
pub fn goldenrod(input string) string { return "\x1b[38;2;216;163;30m${input}\x1b[0m" }
pub fn goldenrod1(input string) string { return "\x1b[38;2;255;191;35m${input}\x1b[0m" }
pub fn goldenrod2(input string) string { return "\x1b[38;2;237;178;33m${input}\x1b[0m" }
pub fn goldenrod3(input string) string { return "\x1b[38;2;204;153;28m${input}\x1b[0m" }
pub fn goldenrod4(input string) string { return "\x1b[38;2;137;104;17m${input}\x1b[0m" }
pub fn floralwhite(input string) string { return "\x1b[38;2;255;249;239m${input}\x1b[0m" }
pub fn darkgoldenrod(input string) string { return "\x1b[38;2;183;132;10m${input}\x1b[0m" }
pub fn darkgoldenrod1(input string) string { return "\x1b[38;2;255;183;12m${input}\x1b[0m" }
pub fn darkgoldenrod2(input string) string { return "\x1b[38;2;237;170;12m${input}\x1b[0m" }
pub fn darkgoldenrod3(input string) string { return "\x1b[38;2;204;147;10m${input}\x1b[0m" }
pub fn darkgoldenrod4(input string) string { return "\x1b[38;2;137;99;7m${input}\x1b[0m" }
pub fn cornsilk(input string) string { return "\x1b[38;2;255;247;219m${input}\x1b[0m" }
pub fn cornsilk2(input string) string { return "\x1b[38;2;237;232;204m${input}\x1b[0m" }
pub fn cornsilk3(input string) string { return "\x1b[38;2;204;198;175m${input}\x1b[0m" }
pub fn lightgoldenrod1(input string) string { return "\x1b[38;2;255;234;137m${input}\x1b[0m" }
pub fn lightgoldenrod2(input string) string { return "\x1b[38;2;237;219;130m${input}\x1b[0m" }
pub fn lightgoldenrod3(input string) string { return "\x1b[38;2;204;188;109m${input}\x1b[0m" }
pub fn gold(input string) string { return "\x1b[38;2;255;214;0m${input}\x1b[0m" }
pub fn gold2(input string) string { return "\x1b[38;2;237;198;0m${input}\x1b[0m" }
pub fn gold3(input string) string { return "\x1b[38;2;204;170;0m${input}\x1b[0m" }
pub fn gold4(input string) string { return "\x1b[38;2;137;114;0m${input}\x1b[0m" }
pub fn cornsilk4(input string) string { return "\x1b[38;2;137;135;119m${input}\x1b[0m" }
pub fn lemonchiffon2(input string) string { return "\x1b[38;2;237;232;188m${input}\x1b[0m" }
pub fn lightgoldenrod(input string) string { return "\x1b[38;2;237;219;130m${input}\x1b[0m" }
pub fn lightgoldenrod4(input string) string { return "\x1b[38;2;137;127;73m${input}\x1b[0m" }
pub fn khaki(input string) string { return "\x1b[38;2;239;229;137m${input}\x1b[0m" }
pub fn khaki1(input string) string { return "\x1b[38;2;255;244;142m${input}\x1b[0m" }
pub fn khaki2(input string) string { return "\x1b[38;2;237;229;132m${input}\x1b[0m" }
pub fn khaki3(input string) string { return "\x1b[38;2;204;196;114m${input}\x1b[0m" }
pub fn khaki4(input string) string { return "\x1b[38;2;137;132;76m${input}\x1b[0m" }
pub fn darkkhaki(input string) string { return "\x1b[38;2;188;181;107m${input}\x1b[0m" }
pub fn lemonchiffon(input string) string { return "\x1b[38;2;255;249;204m${input}\x1b[0m" }
pub fn lemonchiffon3(input string) string { return "\x1b[38;2;204;198;163m${input}\x1b[0m" }
pub fn lemonchiffon4(input string) string { return "\x1b[38;2;137;135;109m${input}\x1b[0m" }
pub fn palegoldenrod(input string) string { return "\x1b[38;2;237;232;168m${input}\x1b[0m" }
pub fn beige(input string) string { return "\x1b[38;2;244;244;219m${input}\x1b[0m" }
pub fn olive(input string) string { return "\x1b[38;2;127;127;0m${input}\x1b[0m" }
pub fn ivory(input string) string { return "\x1b[38;2;255;255;239m${input}\x1b[0m" }
pub fn ivory2(input string) string { return "\x1b[38;2;237;237;221m${input}\x1b[0m" }
pub fn ivory3(input string) string { return "\x1b[38;2;204;204;191m${input}\x1b[0m" }
pub fn ivory4(input string) string { return "\x1b[38;2;137;137;130m${input}\x1b[0m" }
pub fn yellow2(input string) string { return "\x1b[38;2;237;237;0m${input}\x1b[0m" }
pub fn yellow3(input string) string { return "\x1b[38;2;204;204;0m${input}\x1b[0m" }
pub fn yellow4(input string) string { return "\x1b[38;2;137;137;0m${input}\x1b[0m" }
pub fn lightyellow(input string) string { return "\x1b[38;2;255;255;221m${input}\x1b[0m" }
pub fn lightyellow2(input string) string { return "\x1b[38;2;237;237;209m${input}\x1b[0m" }
pub fn lightyellow3(input string) string { return "\x1b[38;2;204;204;178m${input}\x1b[0m" }
pub fn lightyellow4(input string) string { return "\x1b[38;2;137;137;119m${input}\x1b[0m" }
pub fn lightgoldenrodyellow(input string) string { return "\x1b[38;2;249;249;209m${input}\x1b[0m" }
pub fn olivedrab(input string) string { return "\x1b[38;2;107;140;33m${input}\x1b[0m" }
pub fn olivedrab1(input string) string { return "\x1b[38;2;191;255;61m${input}\x1b[0m" }
pub fn olivedrab2(input string) string { return "\x1b[38;2;178;237;56m${input}\x1b[0m" }
pub fn olivedrab3(input string) string { return "\x1b[38;2;153;204;48m${input}\x1b[0m" }
pub fn olivedrab4(input string) string { return "\x1b[38;2;104;137;33m${input}\x1b[0m" }
pub fn darkolivegreen(input string) string { return "\x1b[38;2;84;107;45m${input}\x1b[0m" }
pub fn darkolivegreen1(input string) string { return "\x1b[38;2;201;255;109m${input}\x1b[0m" }
pub fn darkolivegreen2(input string) string { return "\x1b[38;2;186;237;102m${input}\x1b[0m" }
pub fn darkolivegreen3(input string) string { return "\x1b[38;2;160;204;89m${input}\x1b[0m" }
pub fn darkolivegreen4(input string) string { return "\x1b[38;2;109;137;58m${input}\x1b[0m" }
pub fn greenyellow(input string) string { return "\x1b[38;2;170;255;45m${input}\x1b[0m" }
pub fn lawngreen(input string) string { return "\x1b[38;2;122;249;0m${input}\x1b[0m" }
pub fn chartreuse(input string) string { return "\x1b[38;2;124;255;0m${input}\x1b[0m" }
pub fn chartreuse2(input string) string { return "\x1b[38;2;117;237;0m${input}\x1b[0m" }
pub fn chartreuse3(input string) string { return "\x1b[38;2;102;204;0m${input}\x1b[0m" }
pub fn chartreuse4(input string) string { return "\x1b[38;2;68;137;0m${input}\x1b[0m" }
pub fn green2(input string) string { return "\x1b[38;2;0;237;0m${input}\x1b[0m" }
pub fn green3(input string) string { return "\x1b[38;2;0;204;0m${input}\x1b[0m" }
pub fn green4(input string) string { return "\x1b[38;2;0;137;0m${input}\x1b[0m" }
pub fn webgreen(input string) string { return "\x1b[38;2;0;127;0m${input}\x1b[0m" }
pub fn honeydew(input string) string { return "\x1b[38;2;239;255;239m${input}\x1b[0m" }
pub fn honeydew2(input string) string { return "\x1b[38;2;221;237;221m${input}\x1b[0m" }
pub fn honeydew3(input string) string { return "\x1b[38;2;191;204;191m${input}\x1b[0m" }
pub fn honeydew4(input string) string { return "\x1b[38;2;130;137;130m${input}\x1b[0m" }
pub fn darkgreen(input string) string { return "\x1b[38;2;0;99;0m${input}\x1b[0m" }
pub fn palegreen(input string) string { return "\x1b[38;2;150;249;150m${input}\x1b[0m" }
pub fn palegreen1(input string) string { return "\x1b[38;2;153;255;153m${input}\x1b[0m" }
pub fn palegreen3(input string) string { return "\x1b[38;2;122;204;122m${input}\x1b[0m" }
pub fn palegreen4(input string) string { return "\x1b[38;2;81;137;81m${input}\x1b[0m" }
pub fn limegreen(input string) string { return "\x1b[38;2;48;204;48m${input}\x1b[0m" }
pub fn lightgreen(input string) string { return "\x1b[38;2;142;237;142m${input}\x1b[0m" }
pub fn forestgreen(input string) string { return "\x1b[38;2;33;137;33m${input}\x1b[0m" }
pub fn darkseagreen(input string) string { return "\x1b[38;2;142;186;142m${input}\x1b[0m" }
pub fn darkseagreen1(input string) string { return "\x1b[38;2;191;255;191m${input}\x1b[0m" }
pub fn darkseagreen2(input string) string { return "\x1b[38;2;178;237;178m${input}\x1b[0m" }
pub fn darkseagreen3(input string) string { return "\x1b[38;2;153;204;153m${input}\x1b[0m" }
pub fn darkseagreen4(input string) string { return "\x1b[38;2;104;137;104m${input}\x1b[0m" }
pub fn seagreen(input string) string { return "\x1b[38;2;45;137;86m${input}\x1b[0m" }
pub fn seagreen1(input string) string { return "\x1b[38;2;81;255;158m${input}\x1b[0m" }
pub fn seagreen2(input string) string { return "\x1b[38;2;76;237;147m${input}\x1b[0m" }
pub fn seagreen3(input string) string { return "\x1b[38;2;66;204;127m${input}\x1b[0m" }
pub fn mediumseagreen(input string) string { return "\x1b[38;2;58;178;112m${input}\x1b[0m" }
pub fn mintcream(input string) string { return "\x1b[38;2;244;255;249m${input}\x1b[0m" }
pub fn springgreen(input string) string { return "\x1b[38;2;0;255;124m${input}\x1b[0m" }
pub fn springgreen2(input string) string { return "\x1b[38;2;0;237;117m${input}\x1b[0m" }
pub fn springgreen3(input string) string { return "\x1b[38;2;0;204;102m${input}\x1b[0m" }
pub fn springgreen4(input string) string { return "\x1b[38;2;0;137;68m${input}\x1b[0m" }
pub fn mediumspringgreen(input string) string { return "\x1b[38;2;0;249;153m${input}\x1b[0m" }
pub fn aquamarine(input string) string { return "\x1b[38;2;124;255;211m${input}\x1b[0m" }
pub fn aquamarine2(input string) string { return "\x1b[38;2;117;237;196m${input}\x1b[0m" }
pub fn aquamarine3(input string) string { return "\x1b[38;2;102;204;168m${input}\x1b[0m" }
pub fn aquamarine4(input string) string { return "\x1b[38;2;68;137;114m${input}\x1b[0m" }
pub fn turquoise(input string) string { return "\x1b[38;2;63;221;206m${input}\x1b[0m" }
pub fn lightseagreen(input string) string { return "\x1b[38;2;30;175;168m${input}\x1b[0m" }
pub fn mediumturquoise(input string) string { return "\x1b[38;2;71;209;204m${input}\x1b[0m" }
pub fn teal(input string) string { return "\x1b[38;2;0;127;127m${input}\x1b[0m" }
pub fn aqua(input string) string { return "\x1b[38;2;0;255;255m${input}\x1b[0m" }
pub fn cyan2(input string) string { return "\x1b[38;2;0;237;237m${input}\x1b[0m" }
pub fn cyan3(input string) string { return "\x1b[38;2;0;204;204m${input}\x1b[0m" }
pub fn cyan4(input string) string { return "\x1b[38;2;0;137;137m${input}\x1b[0m" }
pub fn azure(input string) string { return "\x1b[38;2;239;255;255m${input}\x1b[0m" }
pub fn azure2(input string) string { return "\x1b[38;2;221;237;237m${input}\x1b[0m" }
pub fn azure3(input string) string { return "\x1b[38;2;191;204;204m${input}\x1b[0m" }
pub fn azure4(input string) string { return "\x1b[38;2;130;137;137m${input}\x1b[0m" }
pub fn cadetblue(input string) string { return "\x1b[38;2;94;158;158m${input}\x1b[0m" }
pub fn lightcyan(input string) string { return "\x1b[38;2;221;255;255m${input}\x1b[0m" }
pub fn lightcyan2(input string) string { return "\x1b[38;2;209;237;237m${input}\x1b[0m" }
pub fn lightcyan3(input string) string { return "\x1b[38;2;178;204;204m${input}\x1b[0m" }
pub fn lightcyan4(input string) string { return "\x1b[38;2;119;137;137m${input}\x1b[0m" }
pub fn turquoise1(input string) string { return "\x1b[38;2;0;244;255m${input}\x1b[0m" }
pub fn turquoise2(input string) string { return "\x1b[38;2;0;226;237m${input}\x1b[0m" }
pub fn turquoise3(input string) string { return "\x1b[38;2;0;196;204m${input}\x1b[0m" }
pub fn turquoise4(input string) string { return "\x1b[38;2;0;132;137m${input}\x1b[0m" }
pub fn darkslategray(input string) string { return "\x1b[38;2;45;79;79m${input}\x1b[0m" }
pub fn darkslategray1(input string) string { return "\x1b[38;2;150;255;255m${input}\x1b[0m" }
pub fn darkslategray2(input string) string { return "\x1b[38;2;140;237;237m${input}\x1b[0m" }
pub fn darkslategray3(input string) string { return "\x1b[38;2;119;204;204m${input}\x1b[0m" }
pub fn darkslategray4(input string) string { return "\x1b[38;2;81;137;137m${input}\x1b[0m" }
pub fn darkturquoise(input string) string { return "\x1b[38;2;0;204;209m${input}\x1b[0m" }
pub fn paleturquoise(input string) string { return "\x1b[38;2;173;237;237m${input}\x1b[0m" }
pub fn paleturquoise1(input string) string { return "\x1b[38;2;186;255;255m${input}\x1b[0m" }
pub fn paleturquoise2(input string) string { return "\x1b[38;2;173;237;237m${input}\x1b[0m" }
pub fn paleturquoise3(input string) string { return "\x1b[38;2;147;204;204m${input}\x1b[0m" }
pub fn paleturquoise4(input string) string { return "\x1b[38;2;102;137;137m${input}\x1b[0m" }
pub fn cadetblue1(input string) string { return "\x1b[38;2;150;244;255m${input}\x1b[0m" }
pub fn cadetblue2(input string) string { return "\x1b[38;2;140;226;237m${input}\x1b[0m" }
pub fn cadetblue3(input string) string { return "\x1b[38;2;119;196;204m${input}\x1b[0m" }
pub fn cadetblue4(input string) string { return "\x1b[38;2;81;132;137m${input}\x1b[0m" }
pub fn powderblue(input string) string { return "\x1b[38;2;175;221;229m${input}\x1b[0m" }
pub fn lightblue4(input string) string { return "\x1b[38;2;102;130;137m${input}\x1b[0m" }
pub fn skyblue(input string) string { return "\x1b[38;2;132;204;234m${input}\x1b[0m" }
pub fn lightblue(input string) string { return "\x1b[38;2;170;214;229m${input}\x1b[0m" }
pub fn lightblue1(input string) string { return "\x1b[38;2;188;237;255m${input}\x1b[0m" }
pub fn lightblue2(input string) string { return "\x1b[38;2;175;221;237m${input}\x1b[0m" }
pub fn lightblue3(input string) string { return "\x1b[38;2;153;191;204m${input}\x1b[0m" }
pub fn deepskyblue(input string) string { return "\x1b[38;2;0;188;255m${input}\x1b[0m" }
pub fn deepskyblue2(input string) string { return "\x1b[38;2;0;175;237m${input}\x1b[0m" }
pub fn deepskyblue3(input string) string { return "\x1b[38;2;0;153;204m${input}\x1b[0m" }
pub fn deepskyblue4(input string) string { return "\x1b[38;2;0;102;137m${input}\x1b[0m" }
pub fn lightskyblue3(input string) string { return "\x1b[38;2;140;181;204m${input}\x1b[0m" }
pub fn skyblue1(input string) string { return "\x1b[38;2;132;204;255m${input}\x1b[0m" }
pub fn skyblue2(input string) string { return "\x1b[38;2;124;191;237m${input}\x1b[0m" }
pub fn skyblue3(input string) string { return "\x1b[38;2;107;165;204m${input}\x1b[0m" }
pub fn skyblue4(input string) string { return "\x1b[38;2;73;109;137m${input}\x1b[0m" }
pub fn lightskyblue(input string) string { return "\x1b[38;2;132;204;249m${input}\x1b[0m" }
pub fn lightskyblue1(input string) string { return "\x1b[38;2;175;224;255m${input}\x1b[0m" }
pub fn lightskyblue2(input string) string { return "\x1b[38;2;163;209;237m${input}\x1b[0m" }
pub fn lightskyblue4(input string) string { return "\x1b[38;2;94;122;137m${input}\x1b[0m" }
pub fn aliceblue(input string) string { return "\x1b[38;2;239;247;255m${input}\x1b[0m" }
pub fn steelblue(input string) string { return "\x1b[38;2;68;130;178m${input}\x1b[0m" }
pub fn steelblue1(input string) string { return "\x1b[38;2;96;183;255m${input}\x1b[0m" }
pub fn steelblue2(input string) string { return "\x1b[38;2;91;170;237m${input}\x1b[0m" }
pub fn steelblue3(input string) string { return "\x1b[38;2;79;147;204m${input}\x1b[0m" }
pub fn steelblue4(input string) string { return "\x1b[38;2;53;99;137m${input}\x1b[0m" }
pub fn slategray(input string) string { return "\x1b[38;2;109;127;142m${input}\x1b[0m" }
pub fn slategray1(input string) string { return "\x1b[38;2;196;224;255m${input}\x1b[0m" }
pub fn slategray2(input string) string { return "\x1b[38;2;183;209;237m${input}\x1b[0m" }
pub fn slategray3(input string) string { return "\x1b[38;2;158;181;204m${input}\x1b[0m" }
pub fn slategray4(input string) string { return "\x1b[38;2;107;122;137m${input}\x1b[0m" }
pub fn dodgerblue(input string) string { return "\x1b[38;2;28;142;255m${input}\x1b[0m" }
pub fn dodgerblue2(input string) string { return "\x1b[38;2;28;132;237m${input}\x1b[0m" }
pub fn dodgerblue3(input string) string { return "\x1b[38;2;22;114;204m${input}\x1b[0m" }
pub fn dodgerblue4(input string) string { return "\x1b[38;2;15;76;137m${input}\x1b[0m" }
pub fn lightslategray(input string) string { return "\x1b[38;2;117;135;153m${input}\x1b[0m" }
pub fn lightsteelblue(input string) string { return "\x1b[38;2;175;193;221m${input}\x1b[0m" }
pub fn lightsteelblue1(input string) string { return "\x1b[38;2;201;224;255m${input}\x1b[0m" }
pub fn lightsteelblue2(input string) string { return "\x1b[38;2;186;209;237m${input}\x1b[0m" }
pub fn lightsteelblue3(input string) string { return "\x1b[38;2;160;181;204m${input}\x1b[0m" }
pub fn lightsteelblue4(input string) string { return "\x1b[38;2;109;122;137m${input}\x1b[0m" }
pub fn cornflowerblue(input string) string { return "\x1b[38;2;99;147;234m${input}\x1b[0m" }
pub fn royalblue(input string) string { return "\x1b[38;2;63;104;224m${input}\x1b[0m" }
pub fn royalblue1(input string) string { return "\x1b[38;2;71;117;255m${input}\x1b[0m" }
pub fn royalblue2(input string) string { return "\x1b[38;2;66;109;237m${input}\x1b[0m" }
pub fn royalblue3(input string) string { return "\x1b[38;2;56;94;204m${input}\x1b[0m" }
pub fn royalblue4(input string) string { return "\x1b[38;2;38;63;137m${input}\x1b[0m" }
pub fn blue2(input string) string { return "\x1b[38;2;0;0;237m${input}\x1b[0m" }
pub fn blue3(input string) string { return "\x1b[38;2;0;0;204m${input}\x1b[0m" }
pub fn blue4(input string) string { return "\x1b[38;2;0;0;137m${input}\x1b[0m" }
pub fn navy(input string) string { return "\x1b[38;2;0;0;127m${input}\x1b[0m" }
pub fn lavender(input string) string { return "\x1b[38;2;229;229;249m${input}\x1b[0m" }
pub fn ghostwhite(input string) string { return "\x1b[38;2;247;247;255m${input}\x1b[0m" }
pub fn midnightblue(input string) string { return "\x1b[38;2;22;22;109m${input}\x1b[0m" }
pub fn slateblue(input string) string { return "\x1b[38;2;104;89;204m${input}\x1b[0m" }
pub fn slateblue1(input string) string { return "\x1b[38;2;130;109;255m${input}\x1b[0m" }
pub fn slateblue3(input string) string { return "\x1b[38;2;104;86;204m${input}\x1b[0m" }
pub fn slateblue4(input string) string { return "\x1b[38;2;68;58;137m${input}\x1b[0m" }
pub fn lightslateblue(input string) string { return "\x1b[38;2;130;109;255m${input}\x1b[0m" }
pub fn slateblue2(input string) string { return "\x1b[38;2;119;102;237m${input}\x1b[0m" }
pub fn darkslateblue(input string) string { return "\x1b[38;2;71;58;137m${input}\x1b[0m" }
pub fn mediumslateblue(input string) string { return "\x1b[38;2;122;102;237m${input}\x1b[0m" }
pub fn mediumpurple(input string) string { return "\x1b[38;2;145;109;216m${input}\x1b[0m" }
pub fn mediumpurple1(input string) string { return "\x1b[38;2;170;130;255m${input}\x1b[0m" }
pub fn mediumpurple2(input string) string { return "\x1b[38;2;158;119;237m${input}\x1b[0m" }
pub fn mediumpurple3(input string) string { return "\x1b[38;2;135;102;204m${input}\x1b[0m" }
pub fn mediumpurple4(input string) string { return "\x1b[38;2;91;68;137m${input}\x1b[0m" }
pub fn purple1(input string) string { return "\x1b[38;2;153;45;255m${input}\x1b[0m" }
pub fn purple2(input string) string { return "\x1b[38;2;142;43;237m${input}\x1b[0m" }
pub fn purple3(input string) string { return "\x1b[38;2;124;35;204m${input}\x1b[0m" }
pub fn purple4(input string) string { return "\x1b[38;2;84;25;137m${input}\x1b[0m" }
pub fn blueviolet(input string) string { return "\x1b[38;2;137;40;224m${input}\x1b[0m" }
pub fn rebeccapurple(input string) string { return "\x1b[38;2;102;51;153m${input}\x1b[0m" }
pub fn indigo(input string) string { return "\x1b[38;2;73;0;130m${input}\x1b[0m" }
pub fn purple(input string) string { return "\x1b[38;2;158;30;239m${input}\x1b[0m" }
pub fn darkorchid(input string) string { return "\x1b[38;2;153;48;204m${input}\x1b[0m" }
pub fn darkorchid1(input string) string { return "\x1b[38;2;188;61;255m${input}\x1b[0m" }
pub fn darkorchid2(input string) string { return "\x1b[38;2;175;56;237m${input}\x1b[0m" }
pub fn darkorchid3(input string) string { return "\x1b[38;2;153;48;204m${input}\x1b[0m" }
pub fn darkorchid4(input string) string { return "\x1b[38;2;102;33;137m${input}\x1b[0m" }
pub fn darkviolet(input string) string { return "\x1b[38;2;147;0;209m${input}\x1b[0m" }
pub fn mediumorchid1(input string) string { return "\x1b[38;2;221;102;255m${input}\x1b[0m" }
pub fn mediumorchid2(input string) string { return "\x1b[38;2;209;94;237m${input}\x1b[0m" }
pub fn mediumorchid3(input string) string { return "\x1b[38;2;178;81;204m${input}\x1b[0m" }
pub fn mediumorchid4(input string) string { return "\x1b[38;2;119;53;137m${input}\x1b[0m" }
pub fn mediumorchid(input string) string { return "\x1b[38;2;183;84;209m${input}\x1b[0m" }
pub fn plum(input string) string { return "\x1b[38;2;219;158;219m${input}\x1b[0m" }
pub fn plum1(input string) string { return "\x1b[38;2;255;186;255m${input}\x1b[0m" }
pub fn plum2(input string) string { return "\x1b[38;2;237;173;237m${input}\x1b[0m" }
pub fn plum3(input string) string { return "\x1b[38;2;204;147;204m${input}\x1b[0m" }
pub fn plum4(input string) string { return "\x1b[38;2;137;102;137m${input}\x1b[0m" }
pub fn orchid(input string) string { return "\x1b[38;2;216;109;211m${input}\x1b[0m" }
pub fn orchid4(input string) string { return "\x1b[38;2;137;68;135m${input}\x1b[0m" }
pub fn violet(input string) string { return "\x1b[38;2;237;130;237m${input}\x1b[0m" }
pub fn magenta2(input string) string { return "\x1b[38;2;237;0;237m${input}\x1b[0m" }
pub fn magenta3(input string) string { return "\x1b[38;2;204;0;204m${input}\x1b[0m" }
pub fn fuchsia(input string) string { return "\x1b[38;2;255;0;255m${input}\x1b[0m" }
pub fn thistle(input string) string { return "\x1b[38;2;214;188;214m${input}\x1b[0m" }
pub fn thistle1(input string) string { return "\x1b[38;2;255;224;255m${input}\x1b[0m" }
pub fn thistle2(input string) string { return "\x1b[38;2;237;209;237m${input}\x1b[0m" }
pub fn thistle3(input string) string { return "\x1b[38;2;204;181;204m${input}\x1b[0m" }
pub fn thistle4(input string) string { return "\x1b[38;2;137;122;137m${input}\x1b[0m" }
pub fn webpurple(input string) string { return "\x1b[38;2;127;0;127m${input}\x1b[0m" }
pub fn darkmagenta(input string) string { return "\x1b[38;2;137;0;137m${input}\x1b[0m" }
pub fn orchid1(input string) string { return "\x1b[38;2;255;130;249m${input}\x1b[0m" }
pub fn orchid2(input string) string { return "\x1b[38;2;237;119;232m${input}\x1b[0m" }
pub fn orchid3(input string) string { return "\x1b[38;2;204;104;198m${input}\x1b[0m" }
pub fn maroon1(input string) string { return "\x1b[38;2;255;51;178m${input}\x1b[0m" }
pub fn maroon2(input string) string { return "\x1b[38;2;237;45;165m${input}\x1b[0m" }
pub fn maroon3(input string) string { return "\x1b[38;2;204;40;142m${input}\x1b[0m" }
pub fn maroon4(input string) string { return "\x1b[38;2;137;28;96m${input}\x1b[0m" }
pub fn violetred(input string) string { return "\x1b[38;2;206;30;142m${input}\x1b[0m" }
pub fn mediumvioletred(input string) string { return "\x1b[38;2;198;20;132m${input}\x1b[0m" }
pub fn deeppink(input string) string { return "\x1b[38;2;255;17;145m${input}\x1b[0m" }
pub fn deeppink2(input string) string { return "\x1b[38;2;237;17;135m${input}\x1b[0m" }
pub fn deeppink4(input string) string { return "\x1b[38;2;137;7;79m${input}\x1b[0m" }
pub fn hotpink(input string) string { return "\x1b[38;2;255;104;178m${input}\x1b[0m" }
pub fn hotpink1(input string) string { return "\x1b[38;2;255;109;178m${input}\x1b[0m" }
pub fn hotpink4(input string) string { return "\x1b[38;2;137;56;96m${input}\x1b[0m" }
pub fn deeppink3(input string) string { return "\x1b[38;2;204;15;117m${input}\x1b[0m" }
pub fn hotpink2(input string) string { return "\x1b[38;2;237;104;165m${input}\x1b[0m" }
pub fn hotpink3(input string) string { return "\x1b[38;2;204;94;142m${input}\x1b[0m" }
pub fn violetred1(input string) string { return "\x1b[38;2;255;61;147m${input}\x1b[0m" }
pub fn violetred2(input string) string { return "\x1b[38;2;237;56;137m${input}\x1b[0m" }
pub fn violetred3(input string) string { return "\x1b[38;2;204;48;119m${input}\x1b[0m" }
pub fn violetred4(input string) string { return "\x1b[38;2;137;33;81m${input}\x1b[0m" }
pub fn maroon(input string) string { return "\x1b[38;2;175;45;94m${input}\x1b[0m" }
pub fn lavenderblush4(input string) string { return "\x1b[38;2;137;130;132m${input}\x1b[0m" }
pub fn lavenderblush(input string) string { return "\x1b[38;2;255;239;244m${input}\x1b[0m" }
pub fn lavenderblush2(input string) string { return "\x1b[38;2;237;221;226m${input}\x1b[0m" }
pub fn lavenderblush3(input string) string { return "\x1b[38;2;204;191;196m${input}\x1b[0m" }
pub fn palevioletred(input string) string { return "\x1b[38;2;216;109;145m${input}\x1b[0m" }
pub fn palevioletred1(input string) string { return "\x1b[38;2;255;130;170m${input}\x1b[0m" }
pub fn palevioletred2(input string) string { return "\x1b[38;2;237;119;158m${input}\x1b[0m" }
pub fn palevioletred3(input string) string { return "\x1b[38;2;204;102;135m${input}\x1b[0m" }
pub fn palevioletred4(input string) string { return "\x1b[38;2;137;68;91m${input}\x1b[0m" }
pub fn pink1(input string) string { return "\x1b[38;2;255;181;196m${input}\x1b[0m" }
pub fn pink2(input string) string { return "\x1b[38;2;237;168;183m${input}\x1b[0m" }
pub fn pink3(input string) string { return "\x1b[38;2;204;142;158m${input}\x1b[0m" }
pub fn pink4(input string) string { return "\x1b[38;2;137;96;107m${input}\x1b[0m" }
pub fn crimson(input string) string { return "\x1b[38;2;219;17;58m${input}\x1b[0m" }
pub fn pink(input string) string { return "\x1b[38;2;255;191;201m${input}\x1b[0m" }
pub fn lightpink(input string) string { return "\x1b[38;2;255;181;191m${input}\x1b[0m" }
pub fn lightpink1(input string) string { return "\x1b[38;2;255;173;183m${input}\x1b[0m" }
pub fn lightpink2(input string) string { return "\x1b[38;2;237;160;170m${input}\x1b[0m" }
pub fn lightpink3(input string) string { return "\x1b[38;2;204;137;147m${input}\x1b[0m" }
pub fn lightpink4(input string) string { return "\x1b[38;2;137;94;99m${input}\x1b[0m" }
pub fn gray1(input string) string { return "\x1b[38;2;2;2;2m${input}\x1b[0m" }
pub fn gray2(input string) string { return "\x1b[38;2;5;5;5m${input}\x1b[0m" }
pub fn gray3(input string) string { return "\x1b[38;2;7;7;7m${input}\x1b[0m" }
pub fn gray4(input string) string { return "\x1b[38;2;7;7;7m${input}\x1b[0m" }
pub fn gray5(input string) string { return "\x1b[38;2;12;12;12m${input}\x1b[0m" }
pub fn gray6(input string) string { return "\x1b[38;2;12;12;12m${input}\x1b[0m" }
pub fn gray7(input string) string { return "\x1b[38;2;17;17;17m${input}\x1b[0m" }
pub fn gray8(input string) string { return "\x1b[38;2;17;17;17m${input}\x1b[0m" }
pub fn gray9(input string) string { return "\x1b[38;2;22;22;22m${input}\x1b[0m" }
pub fn gray10(input string) string { return "\x1b[38;2;25;25;25m${input}\x1b[0m" }
pub fn gray11(input string) string { return "\x1b[38;2;28;28;28m${input}\x1b[0m" }
pub fn gray12(input string) string { return "\x1b[38;2;30;30;30m${input}\x1b[0m" }
pub fn gray13(input string) string { return "\x1b[38;2;30;30;30m${input}\x1b[0m" }
pub fn gray14(input string) string { return "\x1b[38;2;35;35;35m${input}\x1b[0m" }
pub fn gray15(input string) string { return "\x1b[38;2;35;35;35m${input}\x1b[0m" }
pub fn gray16(input string) string { return "\x1b[38;2;40;40;40m${input}\x1b[0m" }
pub fn gray17(input string) string { return "\x1b[38;2;40;40;40m${input}\x1b[0m" }
pub fn gray18(input string) string { return "\x1b[38;2;45;45;45m${input}\x1b[0m" }
pub fn gray19(input string) string { return "\x1b[38;2;45;45;45m${input}\x1b[0m" }
pub fn gray20(input string) string { return "\x1b[38;2;51;51;51m${input}\x1b[0m" }
pub fn gray21(input string) string { return "\x1b[38;2;53;53;53m${input}\x1b[0m" }
pub fn gray22(input string) string { return "\x1b[38;2;56;56;56m${input}\x1b[0m" }
pub fn gray23(input string) string { return "\x1b[38;2;58;58;58m${input}\x1b[0m" }
pub fn gray24(input string) string { return "\x1b[38;2;58;58;58m${input}\x1b[0m" }
pub fn gray25(input string) string { return "\x1b[38;2;63;63;63m${input}\x1b[0m" }
pub fn gray26(input string) string { return "\x1b[38;2;63;63;63m${input}\x1b[0m" }
pub fn gray27(input string) string { return "\x1b[38;2;68;68;68m${input}\x1b[0m" }
pub fn gray28(input string) string { return "\x1b[38;2;68;68;68m${input}\x1b[0m" }
pub fn gray29(input string) string { return "\x1b[38;2;73;73;73m${input}\x1b[0m" }
pub fn gray30(input string) string { return "\x1b[38;2;76;76;76m${input}\x1b[0m" }
pub fn gray31(input string) string { return "\x1b[38;2;79;79;79m${input}\x1b[0m" }
pub fn gray32(input string) string { return "\x1b[38;2;81;81;81m${input}\x1b[0m" }
pub fn gray33(input string) string { return "\x1b[38;2;81;81;81m${input}\x1b[0m" }
pub fn gray34(input string) string { return "\x1b[38;2;86;86;86m${input}\x1b[0m" }
pub fn gray35(input string) string { return "\x1b[38;2;86;86;86m${input}\x1b[0m" }
pub fn gray36(input string) string { return "\x1b[38;2;91;91;91m${input}\x1b[0m" }
pub fn gray37(input string) string { return "\x1b[38;2;91;91;91m${input}\x1b[0m" }
pub fn gray38(input string) string { return "\x1b[38;2;96;96;96m${input}\x1b[0m" }
pub fn gray39(input string) string { return "\x1b[38;2;96;96;96m${input}\x1b[0m" }
pub fn gray40(input string) string { return "\x1b[38;2;102;102;102m${input}\x1b[0m" }
pub fn dimgray(input string) string { return "\x1b[38;2;104;104;104m${input}\x1b[0m" }
pub fn gray42(input string) string { return "\x1b[38;2;107;107;107m${input}\x1b[0m" }
pub fn gray43(input string) string { return "\x1b[38;2;109;109;109m${input}\x1b[0m" }
pub fn gray44(input string) string { return "\x1b[38;2;109;109;109m${input}\x1b[0m" }
pub fn gray45(input string) string { return "\x1b[38;2;114;114;114m${input}\x1b[0m" }
pub fn gray46(input string) string { return "\x1b[38;2;114;114;114m${input}\x1b[0m" }
pub fn gray47(input string) string { return "\x1b[38;2;119;119;119m${input}\x1b[0m" }
pub fn gray48(input string) string { return "\x1b[38;2;119;119;119m${input}\x1b[0m" }
pub fn gray49(input string) string { return "\x1b[38;2;124;124;124m${input}\x1b[0m" }
pub fn gray50(input string) string { return "\x1b[38;2;124;124;124m${input}\x1b[0m" }
pub fn webgray(input string) string { return "\x1b[38;2;127;127;127m${input}\x1b[0m" }
pub fn gray51(input string) string { return "\x1b[38;2;130;130;130m${input}\x1b[0m" }
pub fn gray52(input string) string { return "\x1b[38;2;132;132;132m${input}\x1b[0m" }
pub fn gray53(input string) string { return "\x1b[38;2;132;132;132m${input}\x1b[0m" }
pub fn gray54(input string) string { return "\x1b[38;2;137;137;137m${input}\x1b[0m" }
pub fn gray55(input string) string { return "\x1b[38;2;137;137;137m${input}\x1b[0m" }
pub fn gray56(input string) string { return "\x1b[38;2;142;142;142m${input}\x1b[0m" }
pub fn gray57(input string) string { return "\x1b[38;2;142;142;142m${input}\x1b[0m" }
pub fn gray58(input string) string { return "\x1b[38;2;147;147;147m${input}\x1b[0m" }
pub fn gray59(input string) string { return "\x1b[38;2;147;147;147m${input}\x1b[0m" }
pub fn gray60(input string) string { return "\x1b[38;2;153;153;153m${input}\x1b[0m" }
pub fn gray61(input string) string { return "\x1b[38;2;155;155;155m${input}\x1b[0m" }
pub fn gray62(input string) string { return "\x1b[38;2;158;158;158m${input}\x1b[0m" }
pub fn gray63(input string) string { return "\x1b[38;2;160;160;160m${input}\x1b[0m" }
pub fn gray64(input string) string { return "\x1b[38;2;160;160;160m${input}\x1b[0m" }
pub fn gray65(input string) string { return "\x1b[38;2;165;165;165m${input}\x1b[0m" }
pub fn gray66(input string) string { return "\x1b[38;2;165;165;165m${input}\x1b[0m" }
pub fn darkgray(input string) string { return "\x1b[38;2;168;168;168m${input}\x1b[0m" }
pub fn gray67(input string) string { return "\x1b[38;2;170;170;170m${input}\x1b[0m" }
pub fn gray68(input string) string { return "\x1b[38;2;170;170;170m${input}\x1b[0m" }
pub fn gray69(input string) string { return "\x1b[38;2;175;175;175m${input}\x1b[0m" }
pub fn gray70(input string) string { return "\x1b[38;2;178;178;178m${input}\x1b[0m" }
pub fn gray71(input string) string { return "\x1b[38;2;181;181;181m${input}\x1b[0m" }
pub fn gray72(input string) string { return "\x1b[38;2;183;183;183m${input}\x1b[0m" }
pub fn gray73(input string) string { return "\x1b[38;2;183;183;183m${input}\x1b[0m" }
pub fn gray74(input string) string { return "\x1b[38;2;188;188;188m${input}\x1b[0m" }
pub fn gray(input string) string { return "\x1b[38;2;188;188;188m${input}\x1b[0m" }
pub fn gray75(input string) string { return "\x1b[38;2;188;188;188m${input}\x1b[0m" }
pub fn silver(input string) string { return "\x1b[38;2;191;191;191m${input}\x1b[0m" }
pub fn gray76(input string) string { return "\x1b[38;2;193;193;193m${input}\x1b[0m" }
pub fn gray77(input string) string { return "\x1b[38;2;193;193;193m${input}\x1b[0m" }
pub fn gray78(input string) string { return "\x1b[38;2;198;198;198m${input}\x1b[0m" }
pub fn gray79(input string) string { return "\x1b[38;2;198;198;198m${input}\x1b[0m" }
pub fn gray80(input string) string { return "\x1b[38;2;204;204;204m${input}\x1b[0m" }
pub fn gray81(input string) string { return "\x1b[38;2;206;206;206m${input}\x1b[0m" }
pub fn gray82(input string) string { return "\x1b[38;2;209;209;209m${input}\x1b[0m" }
pub fn lightgray(input string) string { return "\x1b[38;2;209;209;209m${input}\x1b[0m" }
pub fn gray83(input string) string { return "\x1b[38;2;211;211;211m${input}\x1b[0m" }
pub fn gray84(input string) string { return "\x1b[38;2;211;211;211m${input}\x1b[0m" }
pub fn gray85(input string) string { return "\x1b[38;2;216;216;216m${input}\x1b[0m" }
pub fn gray86(input string) string { return "\x1b[38;2;216;216;216m${input}\x1b[0m" }
pub fn gainsboro(input string) string { return "\x1b[38;2;219;219;219m${input}\x1b[0m" }
pub fn gray87(input string) string { return "\x1b[38;2;221;221;221m${input}\x1b[0m" }
pub fn gray88(input string) string { return "\x1b[38;2;221;221;221m${input}\x1b[0m" }
pub fn gray89(input string) string { return "\x1b[38;2;226;226;226m${input}\x1b[0m" }
pub fn gray90(input string) string { return "\x1b[38;2;226;226;226m${input}\x1b[0m" }
pub fn gray91(input string) string { return "\x1b[38;2;232;232;232m${input}\x1b[0m" }
pub fn gray92(input string) string { return "\x1b[38;2;234;234;234m${input}\x1b[0m" }
pub fn gray93(input string) string { return "\x1b[38;2;234;234;234m${input}\x1b[0m" }
pub fn gray94(input string) string { return "\x1b[38;2;239;239;239m${input}\x1b[0m" }
pub fn gray95(input string) string { return "\x1b[38;2;239;239;239m${input}\x1b[0m" }
pub fn gray96(input string) string { return "\x1b[38;2;244;244;244m${input}\x1b[0m" }
pub fn gray97(input string) string { return "\x1b[38;2;244;244;244m${input}\x1b[0m" }
pub fn gray98(input string) string { return "\x1b[38;2;249;249;249m${input}\x1b[0m" }
pub fn gray99(input string) string { return "\x1b[38;2;249;249;249m${input}\x1b[0m" }
pub fn gray100(input string) string { return "\x1b[38;2;255;255;255m${input}\x1b[0m" }

// 256 bit background colour
pub fn on_red2(input string) string { return "\x1b[48;2;237;0;0m${input}\x1b[0m" }
pub fn on_red3(input string) string { return "\x1b[48;2;204;0;0m${input}\x1b[0m" }
pub fn on_snow(input string) string { return "\x1b[48;2;255;249;249m${input}\x1b[0m" }
pub fn on_snow2(input string) string { return "\x1b[48;2;237;232;232m${input}\x1b[0m" }
pub fn on_snow3(input string) string { return "\x1b[48;2;204;198;198m${input}\x1b[0m" }
pub fn on_snow4(input string) string { return "\x1b[48;2;137;135;135m${input}\x1b[0m" }
pub fn on_brown(input string) string { return "\x1b[48;2;163;40;40m${input}\x1b[0m" }
pub fn on_brown1(input string) string { return "\x1b[48;2;255;63;63m${input}\x1b[0m" }
pub fn on_brown2(input string) string { return "\x1b[48;2;237;58;58m${input}\x1b[0m" }
pub fn on_brown3(input string) string { return "\x1b[48;2;204;51;51m${input}\x1b[0m" }
pub fn on_brown4(input string) string { return "\x1b[48;2;137;33;33m${input}\x1b[0m" }
pub fn on_darkred(input string) string { return "\x1b[48;2;137;0;0m${input}\x1b[0m" }
pub fn on_indianred(input string) string { return "\x1b[48;2;204;91;91m${input}\x1b[0m" }
pub fn on_indianred1(input string) string { return "\x1b[48;2;255;104;104m${input}\x1b[0m" }
pub fn on_indianred2(input string) string { return "\x1b[48;2;237;96;96m${input}\x1b[0m" }
pub fn on_indianred3(input string) string { return "\x1b[48;2;204;84;84m${input}\x1b[0m" }
pub fn on_indianred4(input string) string { return "\x1b[48;2;137;56;56m${input}\x1b[0m" }
pub fn on_firebrick(input string) string { return "\x1b[48;2;175;33;33m${input}\x1b[0m" }
pub fn on_firebrick1(input string) string { return "\x1b[48;2;255;45;45m${input}\x1b[0m" }
pub fn on_firebrick2(input string) string { return "\x1b[48;2;237;43;43m${input}\x1b[0m" }
pub fn on_firebrick3(input string) string { return "\x1b[48;2;204;35;35m${input}\x1b[0m" }
pub fn on_firebrick4(input string) string { return "\x1b[48;2;137;25;25m${input}\x1b[0m" }
pub fn on_webmaroon(input string) string { return "\x1b[48;2;127;0;0m${input}\x1b[0m" }
pub fn on_rosybrown(input string) string { return "\x1b[48;2;186;142;142m${input}\x1b[0m" }
pub fn on_rosybrown1(input string) string { return "\x1b[48;2;255;191;191m${input}\x1b[0m" }
pub fn on_rosybrown2(input string) string { return "\x1b[48;2;237;178;178m${input}\x1b[0m" }
pub fn on_rosybrown3(input string) string { return "\x1b[48;2;204;153;153m${input}\x1b[0m" }
pub fn on_rosybrown4(input string) string { return "\x1b[48;2;137;104;104m${input}\x1b[0m" }
pub fn on_lightcoral(input string) string { return "\x1b[48;2;239;127;127m${input}\x1b[0m" }
pub fn on_salmon(input string) string { return "\x1b[48;2;249;127;112m${input}\x1b[0m" }
pub fn on_mistyrose(input string) string { return "\x1b[48;2;255;226;224m${input}\x1b[0m" }
pub fn on_mistyrose2(input string) string { return "\x1b[48;2;237;211;209m${input}\x1b[0m" }
pub fn on_mistyrose3(input string) string { return "\x1b[48;2;204;181;181m${input}\x1b[0m" }
pub fn on_coral1(input string) string { return "\x1b[48;2;255;112;84m${input}\x1b[0m" }
pub fn on_coral2(input string) string { return "\x1b[48;2;237;104;79m${input}\x1b[0m" }
pub fn on_coral3(input string) string { return "\x1b[48;2;204;89;68m${input}\x1b[0m" }
pub fn on_coral4(input string) string { return "\x1b[48;2;137;61;45m${input}\x1b[0m" }
pub fn on_tomato(input string) string { return "\x1b[48;2;255;96;68m${input}\x1b[0m" }
pub fn on_tomato2(input string) string { return "\x1b[48;2;237;91;63m${input}\x1b[0m" }
pub fn on_tomato3(input string) string { return "\x1b[48;2;204;79;56m${input}\x1b[0m" }
pub fn on_tomato4(input string) string { return "\x1b[48;2;137;53;35m${input}\x1b[0m" }
pub fn on_mistyrose4(input string) string { return "\x1b[48;2;137;124;122m${input}\x1b[0m" }
pub fn on_salmon1(input string) string { return "\x1b[48;2;255;137;104m${input}\x1b[0m" }
pub fn on_salmon2(input string) string { return "\x1b[48;2;237;130;96m${input}\x1b[0m" }
pub fn on_salmon3(input string) string { return "\x1b[48;2;204;109;81m${input}\x1b[0m" }
pub fn on_salmon4(input string) string { return "\x1b[48;2;137;73;56m${input}\x1b[0m" }
pub fn on_coral(input string) string { return "\x1b[48;2;255;124;79m${input}\x1b[0m" }
pub fn on_orangered(input string) string { return "\x1b[48;2;255;68;0m${input}\x1b[0m" }
pub fn on_orangered2(input string) string { return "\x1b[48;2;237;63;0m${input}\x1b[0m" }
pub fn on_orangered3(input string) string { return "\x1b[48;2;204;53;0m${input}\x1b[0m" }
pub fn on_orangered4(input string) string { return "\x1b[48;2;137;35;0m${input}\x1b[0m" }
pub fn on_darksalmon(input string) string { return "\x1b[48;2;232;147;119m${input}\x1b[0m" }
pub fn on_lightsalmon(input string) string { return "\x1b[48;2;255;158;119m${input}\x1b[0m" }
pub fn on_lightsalmon2(input string) string { return "\x1b[48;2;237;147;112m${input}\x1b[0m" }
pub fn on_lightsalmon3(input string) string { return "\x1b[48;2;204;127;96m${input}\x1b[0m" }
pub fn on_lightsalmon4(input string) string { return "\x1b[48;2;137;86;63m${input}\x1b[0m" }
pub fn on_sienna(input string) string { return "\x1b[48;2;158;81;43m${input}\x1b[0m" }
pub fn on_sienna1(input string) string { return "\x1b[48;2;255;130;68m${input}\x1b[0m" }
pub fn on_sienna2(input string) string { return "\x1b[48;2;237;119;63m${input}\x1b[0m" }
pub fn on_sienna3(input string) string { return "\x1b[48;2;204;102;56m${input}\x1b[0m" }
pub fn on_sienna4(input string) string { return "\x1b[48;2;137;68;35m${input}\x1b[0m" }
pub fn on_seashell(input string) string { return "\x1b[48;2;255;244;237m${input}\x1b[0m" }
pub fn on_chocolate(input string) string { return "\x1b[48;2;209;104;28m${input}\x1b[0m" }
pub fn on_chocolate1(input string) string { return "\x1b[48;2;255;124;35m${input}\x1b[0m" }
pub fn on_chocolate2(input string) string { return "\x1b[48;2;237;117;30m${input}\x1b[0m" }
pub fn on_chocolate3(input string) string { return "\x1b[48;2;204;102;28m${input}\x1b[0m" }
pub fn on_chocolate4(input string) string { return "\x1b[48;2;137;68;17m${input}\x1b[0m" }
pub fn on_seashell2(input string) string { return "\x1b[48;2;237;226;221m${input}\x1b[0m" }
pub fn on_seashell3(input string) string { return "\x1b[48;2;204;196;188m${input}\x1b[0m" }
pub fn on_seashell4(input string) string { return "\x1b[48;2;137;132;130m${input}\x1b[0m" }
pub fn on_peachpuff(input string) string { return "\x1b[48;2;255;216;183m${input}\x1b[0m" }
pub fn on_peachpuff2(input string) string { return "\x1b[48;2;237;201;170m${input}\x1b[0m" }
pub fn on_peachpuff3(input string) string { return "\x1b[48;2;204;173;147m${input}\x1b[0m" }
pub fn on_peachpuff4(input string) string { return "\x1b[48;2;137;117;99m${input}\x1b[0m" }
pub fn on_sandybrown(input string) string { return "\x1b[48;2;242;163;94m${input}\x1b[0m" }
pub fn on_tan1(input string) string { return "\x1b[48;2;255;163;79m${input}\x1b[0m" }
pub fn on_tan2(input string) string { return "\x1b[48;2;237;153;71m${input}\x1b[0m" }
pub fn on_tan4(input string) string { return "\x1b[48;2;137;89;40m${input}\x1b[0m" }
pub fn on_peru(input string) string { return "\x1b[48;2;204;132;61m${input}\x1b[0m" }
pub fn on_linen(input string) string { return "\x1b[48;2;249;239;229m${input}\x1b[0m" }
pub fn on_bisque3(input string) string { return "\x1b[48;2;204;181;158m${input}\x1b[0m" }
pub fn on_darkorange1(input string) string { return "\x1b[48;2;255;124;0m${input}\x1b[0m" }
pub fn on_darkorange2(input string) string { return "\x1b[48;2;237;117;0m${input}\x1b[0m" }
pub fn on_darkorange3(input string) string { return "\x1b[48;2;204;102;0m${input}\x1b[0m" }
pub fn on_darkorange4(input string) string { return "\x1b[48;2;137;68;0m${input}\x1b[0m" }
pub fn on_tan(input string) string { return "\x1b[48;2;209;178;137m${input}\x1b[0m" }
pub fn on_bisque(input string) string { return "\x1b[48;2;255;226;193m${input}\x1b[0m" }
pub fn on_bisque2(input string) string { return "\x1b[48;2;237;211;181m${input}\x1b[0m" }
pub fn on_bisque4(input string) string { return "\x1b[48;2;137;124;107m${input}\x1b[0m" }
pub fn on_burlywood(input string) string { return "\x1b[48;2;221;183;132m${input}\x1b[0m" }
pub fn on_burlywood1(input string) string { return "\x1b[48;2;255;209;153m${input}\x1b[0m" }
pub fn on_burlywood2(input string) string { return "\x1b[48;2;237;196;142m${input}\x1b[0m" }
pub fn on_burlywood3(input string) string { return "\x1b[48;2;204;168;124m${input}\x1b[0m" }
pub fn on_burlywood4(input string) string { return "\x1b[48;2;137;114;84m${input}\x1b[0m" }
pub fn on_darkorange(input string) string { return "\x1b[48;2;255;137;0m${input}\x1b[0m" }
pub fn on_navajowhite(input string) string { return "\x1b[48;2;255;221;170m${input}\x1b[0m" }
pub fn on_navajowhite2(input string) string { return "\x1b[48;2;237;206;160m${input}\x1b[0m" }
pub fn on_antiquewhite(input string) string { return "\x1b[48;2;249;234;214m${input}\x1b[0m" }
pub fn on_antiquewhite1(input string) string { return "\x1b[48;2;255;237;216m${input}\x1b[0m" }
pub fn on_antiquewhite2(input string) string { return "\x1b[48;2;237;221;204m${input}\x1b[0m" }
pub fn on_antiquewhite3(input string) string { return "\x1b[48;2;204;191;175m${input}\x1b[0m" }
pub fn on_antiquewhite4(input string) string { return "\x1b[48;2;137;130;119m${input}\x1b[0m" }
pub fn on_wheat(input string) string { return "\x1b[48;2;244;221;178m${input}\x1b[0m" }
pub fn on_wheat1(input string) string { return "\x1b[48;2;255;229;183m${input}\x1b[0m" }
pub fn on_wheat2(input string) string { return "\x1b[48;2;237;214;173m${input}\x1b[0m" }
pub fn on_wheat3(input string) string { return "\x1b[48;2;204;183;147m${input}\x1b[0m" }
pub fn on_wheat4(input string) string { return "\x1b[48;2;137;124;102m${input}\x1b[0m" }
pub fn on_orange(input string) string { return "\x1b[48;2;255;163;0m${input}\x1b[0m" }
pub fn on_orange2(input string) string { return "\x1b[48;2;237;153;0m${input}\x1b[0m" }
pub fn on_orange3(input string) string { return "\x1b[48;2;204;132;0m${input}\x1b[0m" }
pub fn on_orange4(input string) string { return "\x1b[48;2;137;89;0m${input}\x1b[0m" }
pub fn on_oldlace(input string) string { return "\x1b[48;2;252;244;229m${input}\x1b[0m" }
pub fn on_moccasin(input string) string { return "\x1b[48;2;255;226;181m${input}\x1b[0m" }
pub fn on_papayawhip(input string) string { return "\x1b[48;2;255;237;211m${input}\x1b[0m" }
pub fn on_navajowhite3(input string) string { return "\x1b[48;2;204;178;137m${input}\x1b[0m" }
pub fn on_navajowhite4(input string) string { return "\x1b[48;2;137;119;91m${input}\x1b[0m" }
pub fn on_blanchedalmond(input string) string { return "\x1b[48;2;255;234;204m${input}\x1b[0m" }
pub fn on_goldenrod(input string) string { return "\x1b[48;2;216;163;30m${input}\x1b[0m" }
pub fn on_goldenrod1(input string) string { return "\x1b[48;2;255;191;35m${input}\x1b[0m" }
pub fn on_goldenrod2(input string) string { return "\x1b[48;2;237;178;33m${input}\x1b[0m" }
pub fn on_goldenrod3(input string) string { return "\x1b[48;2;204;153;28m${input}\x1b[0m" }
pub fn on_goldenrod4(input string) string { return "\x1b[48;2;137;104;17m${input}\x1b[0m" }
pub fn on_floralwhite(input string) string { return "\x1b[48;2;255;249;239m${input}\x1b[0m" }
pub fn on_darkgoldenrod(input string) string { return "\x1b[48;2;183;132;10m${input}\x1b[0m" }
pub fn on_darkgoldenrod1(input string) string { return "\x1b[48;2;255;183;12m${input}\x1b[0m" }
pub fn on_darkgoldenrod2(input string) string { return "\x1b[48;2;237;170;12m${input}\x1b[0m" }
pub fn on_darkgoldenrod3(input string) string { return "\x1b[48;2;204;147;10m${input}\x1b[0m" }
pub fn on_darkgoldenrod4(input string) string { return "\x1b[48;2;137;99;7m${input}\x1b[0m" }
pub fn on_cornsilk(input string) string { return "\x1b[48;2;255;247;219m${input}\x1b[0m" }
pub fn on_cornsilk2(input string) string { return "\x1b[48;2;237;232;204m${input}\x1b[0m" }
pub fn on_cornsilk3(input string) string { return "\x1b[48;2;204;198;175m${input}\x1b[0m" }
pub fn on_lightgoldenrod1(input string) string { return "\x1b[48;2;255;234;137m${input}\x1b[0m" }
pub fn on_lightgoldenrod2(input string) string { return "\x1b[48;2;237;219;130m${input}\x1b[0m" }
pub fn on_lightgoldenrod3(input string) string { return "\x1b[48;2;204;188;109m${input}\x1b[0m" }
pub fn on_gold(input string) string { return "\x1b[48;2;255;214;0m${input}\x1b[0m" }
pub fn on_gold2(input string) string { return "\x1b[48;2;237;198;0m${input}\x1b[0m" }
pub fn on_gold3(input string) string { return "\x1b[48;2;204;170;0m${input}\x1b[0m" }
pub fn on_gold4(input string) string { return "\x1b[48;2;137;114;0m${input}\x1b[0m" }
pub fn on_cornsilk4(input string) string { return "\x1b[48;2;137;135;119m${input}\x1b[0m" }
pub fn on_lemonchiffon2(input string) string { return "\x1b[48;2;237;232;188m${input}\x1b[0m" }
pub fn on_lightgoldenrod(input string) string { return "\x1b[48;2;237;219;130m${input}\x1b[0m" }
pub fn on_lightgoldenrod4(input string) string { return "\x1b[48;2;137;127;73m${input}\x1b[0m" }
pub fn on_khaki(input string) string { return "\x1b[48;2;239;229;137m${input}\x1b[0m" }
pub fn on_khaki1(input string) string { return "\x1b[48;2;255;244;142m${input}\x1b[0m" }
pub fn on_khaki2(input string) string { return "\x1b[48;2;237;229;132m${input}\x1b[0m" }
pub fn on_khaki3(input string) string { return "\x1b[48;2;204;196;114m${input}\x1b[0m" }
pub fn on_khaki4(input string) string { return "\x1b[48;2;137;132;76m${input}\x1b[0m" }
pub fn on_darkkhaki(input string) string { return "\x1b[48;2;188;181;107m${input}\x1b[0m" }
pub fn on_lemonchiffon(input string) string { return "\x1b[48;2;255;249;204m${input}\x1b[0m" }
pub fn on_lemonchiffon3(input string) string { return "\x1b[48;2;204;198;163m${input}\x1b[0m" }
pub fn on_lemonchiffon4(input string) string { return "\x1b[48;2;137;135;109m${input}\x1b[0m" }
pub fn on_palegoldenrod(input string) string { return "\x1b[48;2;237;232;168m${input}\x1b[0m" }
pub fn on_beige(input string) string { return "\x1b[48;2;244;244;219m${input}\x1b[0m" }
pub fn on_olive(input string) string { return "\x1b[48;2;127;127;0m${input}\x1b[0m" }
pub fn on_ivory(input string) string { return "\x1b[48;2;255;255;239m${input}\x1b[0m" }
pub fn on_ivory2(input string) string { return "\x1b[48;2;237;237;221m${input}\x1b[0m" }
pub fn on_ivory3(input string) string { return "\x1b[48;2;204;204;191m${input}\x1b[0m" }
pub fn on_ivory4(input string) string { return "\x1b[48;2;137;137;130m${input}\x1b[0m" }
pub fn on_yellow2(input string) string { return "\x1b[48;2;237;237;0m${input}\x1b[0m" }
pub fn on_yellow3(input string) string { return "\x1b[48;2;204;204;0m${input}\x1b[0m" }
pub fn on_yellow4(input string) string { return "\x1b[48;2;137;137;0m${input}\x1b[0m" }
pub fn on_lightyellow(input string) string { return "\x1b[48;2;255;255;221m${input}\x1b[0m" }
pub fn on_lightyellow2(input string) string { return "\x1b[48;2;237;237;209m${input}\x1b[0m" }
pub fn on_lightyellow3(input string) string { return "\x1b[48;2;204;204;178m${input}\x1b[0m" }
pub fn on_lightyellow4(input string) string { return "\x1b[48;2;137;137;119m${input}\x1b[0m" }
pub fn on_lightgoldenrodyellow(input string) string { return "\x1b[48;2;249;249;209m${input}\x1b[0m" }
pub fn on_olivedrab(input string) string { return "\x1b[48;2;107;140;33m${input}\x1b[0m" }
pub fn on_olivedrab1(input string) string { return "\x1b[48;2;191;255;61m${input}\x1b[0m" }
pub fn on_olivedrab2(input string) string { return "\x1b[48;2;178;237;56m${input}\x1b[0m" }
pub fn on_olivedrab3(input string) string { return "\x1b[48;2;153;204;48m${input}\x1b[0m" }
pub fn on_olivedrab4(input string) string { return "\x1b[48;2;104;137;33m${input}\x1b[0m" }
pub fn on_darkolivegreen(input string) string { return "\x1b[48;2;84;107;45m${input}\x1b[0m" }
pub fn on_darkolivegreen1(input string) string { return "\x1b[48;2;201;255;109m${input}\x1b[0m" }
pub fn on_darkolivegreen2(input string) string { return "\x1b[48;2;186;237;102m${input}\x1b[0m" }
pub fn on_darkolivegreen3(input string) string { return "\x1b[48;2;160;204;89m${input}\x1b[0m" }
pub fn on_darkolivegreen4(input string) string { return "\x1b[48;2;109;137;58m${input}\x1b[0m" }
pub fn on_greenyellow(input string) string { return "\x1b[48;2;170;255;45m${input}\x1b[0m" }
pub fn on_lawngreen(input string) string { return "\x1b[48;2;122;249;0m${input}\x1b[0m" }
pub fn on_chartreuse(input string) string { return "\x1b[48;2;124;255;0m${input}\x1b[0m" }
pub fn on_chartreuse2(input string) string { return "\x1b[48;2;117;237;0m${input}\x1b[0m" }
pub fn on_chartreuse3(input string) string { return "\x1b[48;2;102;204;0m${input}\x1b[0m" }
pub fn on_chartreuse4(input string) string { return "\x1b[48;2;68;137;0m${input}\x1b[0m" }
pub fn on_green2(input string) string { return "\x1b[48;2;0;237;0m${input}\x1b[0m" }
pub fn on_green3(input string) string { return "\x1b[48;2;0;204;0m${input}\x1b[0m" }
pub fn on_green4(input string) string { return "\x1b[48;2;0;137;0m${input}\x1b[0m" }
pub fn on_webgreen(input string) string { return "\x1b[48;2;0;127;0m${input}\x1b[0m" }
pub fn on_honeydew(input string) string { return "\x1b[48;2;239;255;239m${input}\x1b[0m" }
pub fn on_honeydew2(input string) string { return "\x1b[48;2;221;237;221m${input}\x1b[0m" }
pub fn on_honeydew3(input string) string { return "\x1b[48;2;191;204;191m${input}\x1b[0m" }
pub fn on_honeydew4(input string) string { return "\x1b[48;2;130;137;130m${input}\x1b[0m" }
pub fn on_darkgreen(input string) string { return "\x1b[48;2;0;99;0m${input}\x1b[0m" }
pub fn on_palegreen(input string) string { return "\x1b[48;2;150;249;150m${input}\x1b[0m" }
pub fn on_palegreen1(input string) string { return "\x1b[48;2;153;255;153m${input}\x1b[0m" }
pub fn on_palegreen3(input string) string { return "\x1b[48;2;122;204;122m${input}\x1b[0m" }
pub fn on_palegreen4(input string) string { return "\x1b[48;2;81;137;81m${input}\x1b[0m" }
pub fn on_limegreen(input string) string { return "\x1b[48;2;48;204;48m${input}\x1b[0m" }
pub fn on_lightgreen(input string) string { return "\x1b[48;2;142;237;142m${input}\x1b[0m" }
pub fn on_forestgreen(input string) string { return "\x1b[48;2;33;137;33m${input}\x1b[0m" }
pub fn on_darkseagreen(input string) string { return "\x1b[48;2;142;186;142m${input}\x1b[0m" }
pub fn on_darkseagreen1(input string) string { return "\x1b[48;2;191;255;191m${input}\x1b[0m" }
pub fn on_darkseagreen2(input string) string { return "\x1b[48;2;178;237;178m${input}\x1b[0m" }
pub fn on_darkseagreen3(input string) string { return "\x1b[48;2;153;204;153m${input}\x1b[0m" }
pub fn on_darkseagreen4(input string) string { return "\x1b[48;2;104;137;104m${input}\x1b[0m" }
pub fn on_seagreen(input string) string { return "\x1b[48;2;45;137;86m${input}\x1b[0m" }
pub fn on_seagreen1(input string) string { return "\x1b[48;2;81;255;158m${input}\x1b[0m" }
pub fn on_seagreen2(input string) string { return "\x1b[48;2;76;237;147m${input}\x1b[0m" }
pub fn on_seagreen3(input string) string { return "\x1b[48;2;66;204;127m${input}\x1b[0m" }
pub fn on_mediumseagreen(input string) string { return "\x1b[48;2;58;178;112m${input}\x1b[0m" }
pub fn on_mintcream(input string) string { return "\x1b[48;2;244;255;249m${input}\x1b[0m" }
pub fn on_springgreen(input string) string { return "\x1b[48;2;0;255;124m${input}\x1b[0m" }
pub fn on_springgreen2(input string) string { return "\x1b[48;2;0;237;117m${input}\x1b[0m" }
pub fn on_springgreen3(input string) string { return "\x1b[48;2;0;204;102m${input}\x1b[0m" }
pub fn on_springgreen4(input string) string { return "\x1b[48;2;0;137;68m${input}\x1b[0m" }
pub fn on_mediumspringgreen(input string) string { return "\x1b[48;2;0;249;153m${input}\x1b[0m" }
pub fn on_aquamarine(input string) string { return "\x1b[48;2;124;255;211m${input}\x1b[0m" }
pub fn on_aquamarine2(input string) string { return "\x1b[48;2;117;237;196m${input}\x1b[0m" }
pub fn on_aquamarine3(input string) string { return "\x1b[48;2;102;204;168m${input}\x1b[0m" }
pub fn on_aquamarine4(input string) string { return "\x1b[48;2;68;137;114m${input}\x1b[0m" }
pub fn on_turquoise(input string) string { return "\x1b[48;2;63;221;206m${input}\x1b[0m" }
pub fn on_lightseagreen(input string) string { return "\x1b[48;2;30;175;168m${input}\x1b[0m" }
pub fn on_mediumturquoise(input string) string { return "\x1b[48;2;71;209;204m${input}\x1b[0m" }
pub fn on_teal(input string) string { return "\x1b[48;2;0;127;127m${input}\x1b[0m" }
pub fn on_aqua(input string) string { return "\x1b[48;2;0;255;255m${input}\x1b[0m" }
pub fn on_cyan2(input string) string { return "\x1b[48;2;0;237;237m${input}\x1b[0m" }
pub fn on_cyan3(input string) string { return "\x1b[48;2;0;204;204m${input}\x1b[0m" }
pub fn on_cyan4(input string) string { return "\x1b[48;2;0;137;137m${input}\x1b[0m" }
pub fn on_azure(input string) string { return "\x1b[48;2;239;255;255m${input}\x1b[0m" }
pub fn on_azure2(input string) string { return "\x1b[48;2;221;237;237m${input}\x1b[0m" }
pub fn on_azure3(input string) string { return "\x1b[48;2;191;204;204m${input}\x1b[0m" }
pub fn on_azure4(input string) string { return "\x1b[48;2;130;137;137m${input}\x1b[0m" }
pub fn on_cadetblue(input string) string { return "\x1b[48;2;94;158;158m${input}\x1b[0m" }
pub fn on_lightcyan(input string) string { return "\x1b[48;2;221;255;255m${input}\x1b[0m" }
pub fn on_lightcyan2(input string) string { return "\x1b[48;2;209;237;237m${input}\x1b[0m" }
pub fn on_lightcyan3(input string) string { return "\x1b[48;2;178;204;204m${input}\x1b[0m" }
pub fn on_lightcyan4(input string) string { return "\x1b[48;2;119;137;137m${input}\x1b[0m" }
pub fn on_turquoise1(input string) string { return "\x1b[48;2;0;244;255m${input}\x1b[0m" }
pub fn on_turquoise2(input string) string { return "\x1b[48;2;0;226;237m${input}\x1b[0m" }
pub fn on_turquoise3(input string) string { return "\x1b[48;2;0;196;204m${input}\x1b[0m" }
pub fn on_turquoise4(input string) string { return "\x1b[48;2;0;132;137m${input}\x1b[0m" }
pub fn on_darkslategray(input string) string { return "\x1b[48;2;45;79;79m${input}\x1b[0m" }
pub fn on_darkslategray1(input string) string { return "\x1b[48;2;150;255;255m${input}\x1b[0m" }
pub fn on_darkslategray2(input string) string { return "\x1b[48;2;140;237;237m${input}\x1b[0m" }
pub fn on_darkslategray3(input string) string { return "\x1b[48;2;119;204;204m${input}\x1b[0m" }
pub fn on_darkslategray4(input string) string { return "\x1b[48;2;81;137;137m${input}\x1b[0m" }
pub fn on_darkturquoise(input string) string { return "\x1b[48;2;0;204;209m${input}\x1b[0m" }
pub fn on_paleturquoise(input string) string { return "\x1b[48;2;173;237;237m${input}\x1b[0m" }
pub fn on_paleturquoise1(input string) string { return "\x1b[48;2;186;255;255m${input}\x1b[0m" }
pub fn on_paleturquoise2(input string) string { return "\x1b[48;2;173;237;237m${input}\x1b[0m" }
pub fn on_paleturquoise3(input string) string { return "\x1b[48;2;147;204;204m${input}\x1b[0m" }
pub fn on_paleturquoise4(input string) string { return "\x1b[48;2;102;137;137m${input}\x1b[0m" }
pub fn on_cadetblue1(input string) string { return "\x1b[48;2;150;244;255m${input}\x1b[0m" }
pub fn on_cadetblue2(input string) string { return "\x1b[48;2;140;226;237m${input}\x1b[0m" }
pub fn on_cadetblue3(input string) string { return "\x1b[48;2;119;196;204m${input}\x1b[0m" }
pub fn on_cadetblue4(input string) string { return "\x1b[48;2;81;132;137m${input}\x1b[0m" }
pub fn on_powderblue(input string) string { return "\x1b[48;2;175;221;229m${input}\x1b[0m" }
pub fn on_lightblue4(input string) string { return "\x1b[48;2;102;130;137m${input}\x1b[0m" }
pub fn on_skyblue(input string) string { return "\x1b[48;2;132;204;234m${input}\x1b[0m" }
pub fn on_lightblue(input string) string { return "\x1b[48;2;170;214;229m${input}\x1b[0m" }
pub fn on_lightblue1(input string) string { return "\x1b[48;2;188;237;255m${input}\x1b[0m" }
pub fn on_lightblue2(input string) string { return "\x1b[48;2;175;221;237m${input}\x1b[0m" }
pub fn on_lightblue3(input string) string { return "\x1b[48;2;153;191;204m${input}\x1b[0m" }
pub fn on_deepskyblue(input string) string { return "\x1b[48;2;0;188;255m${input}\x1b[0m" }
pub fn on_deepskyblue2(input string) string { return "\x1b[48;2;0;175;237m${input}\x1b[0m" }
pub fn on_deepskyblue3(input string) string { return "\x1b[48;2;0;153;204m${input}\x1b[0m" }
pub fn on_deepskyblue4(input string) string { return "\x1b[48;2;0;102;137m${input}\x1b[0m" }
pub fn on_lightskyblue3(input string) string { return "\x1b[48;2;140;181;204m${input}\x1b[0m" }
pub fn on_skyblue1(input string) string { return "\x1b[48;2;132;204;255m${input}\x1b[0m" }
pub fn on_skyblue2(input string) string { return "\x1b[48;2;124;191;237m${input}\x1b[0m" }
pub fn on_skyblue3(input string) string { return "\x1b[48;2;107;165;204m${input}\x1b[0m" }
pub fn on_skyblue4(input string) string { return "\x1b[48;2;73;109;137m${input}\x1b[0m" }
pub fn on_lightskyblue(input string) string { return "\x1b[48;2;132;204;249m${input}\x1b[0m" }
pub fn on_lightskyblue1(input string) string { return "\x1b[48;2;175;224;255m${input}\x1b[0m" }
pub fn on_lightskyblue2(input string) string { return "\x1b[48;2;163;209;237m${input}\x1b[0m" }
pub fn on_lightskyblue4(input string) string { return "\x1b[48;2;94;122;137m${input}\x1b[0m" }
pub fn on_aliceblue(input string) string { return "\x1b[48;2;239;247;255m${input}\x1b[0m" }
pub fn on_steelblue(input string) string { return "\x1b[48;2;68;130;178m${input}\x1b[0m" }
pub fn on_steelblue1(input string) string { return "\x1b[48;2;96;183;255m${input}\x1b[0m" }
pub fn on_steelblue2(input string) string { return "\x1b[48;2;91;170;237m${input}\x1b[0m" }
pub fn on_steelblue3(input string) string { return "\x1b[48;2;79;147;204m${input}\x1b[0m" }
pub fn on_steelblue4(input string) string { return "\x1b[48;2;53;99;137m${input}\x1b[0m" }
pub fn on_slategray(input string) string { return "\x1b[48;2;109;127;142m${input}\x1b[0m" }
pub fn on_slategray1(input string) string { return "\x1b[48;2;196;224;255m${input}\x1b[0m" }
pub fn on_slategray2(input string) string { return "\x1b[48;2;183;209;237m${input}\x1b[0m" }
pub fn on_slategray3(input string) string { return "\x1b[48;2;158;181;204m${input}\x1b[0m" }
pub fn on_slategray4(input string) string { return "\x1b[48;2;107;122;137m${input}\x1b[0m" }
pub fn on_dodgerblue(input string) string { return "\x1b[48;2;28;142;255m${input}\x1b[0m" }
pub fn on_dodgerblue2(input string) string { return "\x1b[48;2;28;132;237m${input}\x1b[0m" }
pub fn on_dodgerblue3(input string) string { return "\x1b[48;2;22;114;204m${input}\x1b[0m" }
pub fn on_dodgerblue4(input string) string { return "\x1b[48;2;15;76;137m${input}\x1b[0m" }
pub fn on_lightslategray(input string) string { return "\x1b[48;2;117;135;153m${input}\x1b[0m" }
pub fn on_lightsteelblue(input string) string { return "\x1b[48;2;175;193;221m${input}\x1b[0m" }
pub fn on_lightsteelblue1(input string) string { return "\x1b[48;2;201;224;255m${input}\x1b[0m" }
pub fn on_lightsteelblue2(input string) string { return "\x1b[48;2;186;209;237m${input}\x1b[0m" }
pub fn on_lightsteelblue3(input string) string { return "\x1b[48;2;160;181;204m${input}\x1b[0m" }
pub fn on_lightsteelblue4(input string) string { return "\x1b[48;2;109;122;137m${input}\x1b[0m" }
pub fn on_cornflowerblue(input string) string { return "\x1b[48;2;99;147;234m${input}\x1b[0m" }
pub fn on_royalblue(input string) string { return "\x1b[48;2;63;104;224m${input}\x1b[0m" }
pub fn on_royalblue1(input string) string { return "\x1b[48;2;71;117;255m${input}\x1b[0m" }
pub fn on_royalblue2(input string) string { return "\x1b[48;2;66;109;237m${input}\x1b[0m" }
pub fn on_royalblue3(input string) string { return "\x1b[48;2;56;94;204m${input}\x1b[0m" }
pub fn on_royalblue4(input string) string { return "\x1b[48;2;38;63;137m${input}\x1b[0m" }
pub fn on_blue2(input string) string { return "\x1b[48;2;0;0;237m${input}\x1b[0m" }
pub fn on_blue3(input string) string { return "\x1b[48;2;0;0;204m${input}\x1b[0m" }
pub fn on_blue4(input string) string { return "\x1b[48;2;0;0;137m${input}\x1b[0m" }
pub fn on_navy(input string) string { return "\x1b[48;2;0;0;127m${input}\x1b[0m" }
pub fn on_lavender(input string) string { return "\x1b[48;2;229;229;249m${input}\x1b[0m" }
pub fn on_ghostwhite(input string) string { return "\x1b[48;2;247;247;255m${input}\x1b[0m" }
pub fn on_midnightblue(input string) string { return "\x1b[48;2;22;22;109m${input}\x1b[0m" }
pub fn on_slateblue(input string) string { return "\x1b[48;2;104;89;204m${input}\x1b[0m" }
pub fn on_slateblue1(input string) string { return "\x1b[48;2;130;109;255m${input}\x1b[0m" }
pub fn on_slateblue3(input string) string { return "\x1b[48;2;104;86;204m${input}\x1b[0m" }
pub fn on_slateblue4(input string) string { return "\x1b[48;2;68;58;137m${input}\x1b[0m" }
pub fn on_lightslateblue(input string) string { return "\x1b[48;2;130;109;255m${input}\x1b[0m" }
pub fn on_slateblue2(input string) string { return "\x1b[48;2;119;102;237m${input}\x1b[0m" }
pub fn on_darkslateblue(input string) string { return "\x1b[48;2;71;58;137m${input}\x1b[0m" }
pub fn on_mediumslateblue(input string) string { return "\x1b[48;2;122;102;237m${input}\x1b[0m" }
pub fn on_mediumpurple(input string) string { return "\x1b[48;2;145;109;216m${input}\x1b[0m" }
pub fn on_mediumpurple1(input string) string { return "\x1b[48;2;170;130;255m${input}\x1b[0m" }
pub fn on_mediumpurple2(input string) string { return "\x1b[48;2;158;119;237m${input}\x1b[0m" }
pub fn on_mediumpurple3(input string) string { return "\x1b[48;2;135;102;204m${input}\x1b[0m" }
pub fn on_mediumpurple4(input string) string { return "\x1b[48;2;91;68;137m${input}\x1b[0m" }
pub fn on_purple1(input string) string { return "\x1b[48;2;153;45;255m${input}\x1b[0m" }
pub fn on_purple2(input string) string { return "\x1b[48;2;142;43;237m${input}\x1b[0m" }
pub fn on_purple3(input string) string { return "\x1b[48;2;124;35;204m${input}\x1b[0m" }
pub fn on_purple4(input string) string { return "\x1b[48;2;84;25;137m${input}\x1b[0m" }
pub fn on_blueviolet(input string) string { return "\x1b[48;2;137;40;224m${input}\x1b[0m" }
pub fn on_rebeccapurple(input string) string { return "\x1b[48;2;102;51;153m${input}\x1b[0m" }
pub fn on_indigo(input string) string { return "\x1b[48;2;73;0;130m${input}\x1b[0m" }
pub fn on_purple(input string) string { return "\x1b[48;2;158;30;239m${input}\x1b[0m" }
pub fn on_darkorchid(input string) string { return "\x1b[48;2;153;48;204m${input}\x1b[0m" }
pub fn on_darkorchid1(input string) string { return "\x1b[48;2;188;61;255m${input}\x1b[0m" }
pub fn on_darkorchid2(input string) string { return "\x1b[48;2;175;56;237m${input}\x1b[0m" }
pub fn on_darkorchid3(input string) string { return "\x1b[48;2;153;48;204m${input}\x1b[0m" }
pub fn on_darkorchid4(input string) string { return "\x1b[48;2;102;33;137m${input}\x1b[0m" }
pub fn on_darkviolet(input string) string { return "\x1b[48;2;147;0;209m${input}\x1b[0m" }
pub fn on_mediumorchid1(input string) string { return "\x1b[48;2;221;102;255m${input}\x1b[0m" }
pub fn on_mediumorchid2(input string) string { return "\x1b[48;2;209;94;237m${input}\x1b[0m" }
pub fn on_mediumorchid3(input string) string { return "\x1b[48;2;178;81;204m${input}\x1b[0m" }
pub fn on_mediumorchid4(input string) string { return "\x1b[48;2;119;53;137m${input}\x1b[0m" }
pub fn on_mediumorchid(input string) string { return "\x1b[48;2;183;84;209m${input}\x1b[0m" }
pub fn on_plum(input string) string { return "\x1b[48;2;219;158;219m${input}\x1b[0m" }
pub fn on_plum1(input string) string { return "\x1b[48;2;255;186;255m${input}\x1b[0m" }
pub fn on_plum2(input string) string { return "\x1b[48;2;237;173;237m${input}\x1b[0m" }
pub fn on_plum3(input string) string { return "\x1b[48;2;204;147;204m${input}\x1b[0m" }
pub fn on_plum4(input string) string { return "\x1b[48;2;137;102;137m${input}\x1b[0m" }
pub fn on_orchid(input string) string { return "\x1b[48;2;216;109;211m${input}\x1b[0m" }
pub fn on_orchid4(input string) string { return "\x1b[48;2;137;68;135m${input}\x1b[0m" }
pub fn on_violet(input string) string { return "\x1b[48;2;237;130;237m${input}\x1b[0m" }
pub fn on_magenta2(input string) string { return "\x1b[48;2;237;0;237m${input}\x1b[0m" }
pub fn on_magenta3(input string) string { return "\x1b[48;2;204;0;204m${input}\x1b[0m" }
pub fn on_fuchsia(input string) string { return "\x1b[48;2;255;0;255m${input}\x1b[0m" }
pub fn on_thistle(input string) string { return "\x1b[48;2;214;188;214m${input}\x1b[0m" }
pub fn on_thistle1(input string) string { return "\x1b[48;2;255;224;255m${input}\x1b[0m" }
pub fn on_thistle2(input string) string { return "\x1b[48;2;237;209;237m${input}\x1b[0m" }
pub fn on_thistle3(input string) string { return "\x1b[48;2;204;181;204m${input}\x1b[0m" }
pub fn on_thistle4(input string) string { return "\x1b[48;2;137;122;137m${input}\x1b[0m" }
pub fn on_webpurple(input string) string { return "\x1b[48;2;127;0;127m${input}\x1b[0m" }
pub fn on_darkmagenta(input string) string { return "\x1b[48;2;137;0;137m${input}\x1b[0m" }
pub fn on_orchid1(input string) string { return "\x1b[48;2;255;130;249m${input}\x1b[0m" }
pub fn on_orchid2(input string) string { return "\x1b[48;2;237;119;232m${input}\x1b[0m" }
pub fn on_orchid3(input string) string { return "\x1b[48;2;204;104;198m${input}\x1b[0m" }
pub fn on_maroon1(input string) string { return "\x1b[48;2;255;51;178m${input}\x1b[0m" }
pub fn on_maroon2(input string) string { return "\x1b[48;2;237;45;165m${input}\x1b[0m" }
pub fn on_maroon3(input string) string { return "\x1b[48;2;204;40;142m${input}\x1b[0m" }
pub fn on_maroon4(input string) string { return "\x1b[48;2;137;28;96m${input}\x1b[0m" }
pub fn on_violetred(input string) string { return "\x1b[48;2;206;30;142m${input}\x1b[0m" }
pub fn on_mediumvioletred(input string) string { return "\x1b[48;2;198;20;132m${input}\x1b[0m" }
pub fn on_deeppink(input string) string { return "\x1b[48;2;255;17;145m${input}\x1b[0m" }
pub fn on_deeppink2(input string) string { return "\x1b[48;2;237;17;135m${input}\x1b[0m" }
pub fn on_deeppink4(input string) string { return "\x1b[48;2;137;7;79m${input}\x1b[0m" }
pub fn on_hotpink(input string) string { return "\x1b[48;2;255;104;178m${input}\x1b[0m" }
pub fn on_hotpink1(input string) string { return "\x1b[48;2;255;109;178m${input}\x1b[0m" }
pub fn on_hotpink4(input string) string { return "\x1b[48;2;137;56;96m${input}\x1b[0m" }
pub fn on_deeppink3(input string) string { return "\x1b[48;2;204;15;117m${input}\x1b[0m" }
pub fn on_hotpink2(input string) string { return "\x1b[48;2;237;104;165m${input}\x1b[0m" }
pub fn on_hotpink3(input string) string { return "\x1b[48;2;204;94;142m${input}\x1b[0m" }
pub fn on_violetred1(input string) string { return "\x1b[48;2;255;61;147m${input}\x1b[0m" }
pub fn on_violetred2(input string) string { return "\x1b[48;2;237;56;137m${input}\x1b[0m" }
pub fn on_violetred3(input string) string { return "\x1b[48;2;204;48;119m${input}\x1b[0m" }
pub fn on_violetred4(input string) string { return "\x1b[48;2;137;33;81m${input}\x1b[0m" }
pub fn on_maroon(input string) string { return "\x1b[48;2;175;45;94m${input}\x1b[0m" }
pub fn on_lavenderblush4(input string) string { return "\x1b[48;2;137;130;132m${input}\x1b[0m" }
pub fn on_lavenderblush(input string) string { return "\x1b[48;2;255;239;244m${input}\x1b[0m" }
pub fn on_lavenderblush2(input string) string { return "\x1b[48;2;237;221;226m${input}\x1b[0m" }
pub fn on_lavenderblush3(input string) string { return "\x1b[48;2;204;191;196m${input}\x1b[0m" }
pub fn on_palevioletred(input string) string { return "\x1b[48;2;216;109;145m${input}\x1b[0m" }
pub fn on_palevioletred1(input string) string { return "\x1b[48;2;255;130;170m${input}\x1b[0m" }
pub fn on_palevioletred2(input string) string { return "\x1b[48;2;237;119;158m${input}\x1b[0m" }
pub fn on_palevioletred3(input string) string { return "\x1b[48;2;204;102;135m${input}\x1b[0m" }
pub fn on_palevioletred4(input string) string { return "\x1b[48;2;137;68;91m${input}\x1b[0m" }
pub fn on_pink1(input string) string { return "\x1b[48;2;255;181;196m${input}\x1b[0m" }
pub fn on_pink2(input string) string { return "\x1b[48;2;237;168;183m${input}\x1b[0m" }
pub fn on_pink3(input string) string { return "\x1b[48;2;204;142;158m${input}\x1b[0m" }
pub fn on_pink4(input string) string { return "\x1b[48;2;137;96;107m${input}\x1b[0m" }
pub fn on_crimson(input string) string { return "\x1b[48;2;219;17;58m${input}\x1b[0m" }
pub fn on_pink(input string) string { return "\x1b[48;2;255;191;201m${input}\x1b[0m" }
pub fn on_lightpink(input string) string { return "\x1b[48;2;255;181;191m${input}\x1b[0m" }
pub fn on_lightpink1(input string) string { return "\x1b[48;2;255;173;183m${input}\x1b[0m" }
pub fn on_lightpink2(input string) string { return "\x1b[48;2;237;160;170m${input}\x1b[0m" }
pub fn on_lightpink3(input string) string { return "\x1b[48;2;204;137;147m${input}\x1b[0m" }
pub fn on_lightpink4(input string) string { return "\x1b[48;2;137;94;99m${input}\x1b[0m" }
pub fn on_gray1(input string) string { return "\x1b[48;2;2;2;2m${input}\x1b[0m" }
pub fn on_gray2(input string) string { return "\x1b[48;2;5;5;5m${input}\x1b[0m" }
pub fn on_gray3(input string) string { return "\x1b[48;2;7;7;7m${input}\x1b[0m" }
pub fn on_gray4(input string) string { return "\x1b[48;2;7;7;7m${input}\x1b[0m" }
pub fn on_gray5(input string) string { return "\x1b[48;2;12;12;12m${input}\x1b[0m" }
pub fn on_gray6(input string) string { return "\x1b[48;2;12;12;12m${input}\x1b[0m" }
pub fn on_gray7(input string) string { return "\x1b[48;2;17;17;17m${input}\x1b[0m" }
pub fn on_gray8(input string) string { return "\x1b[48;2;17;17;17m${input}\x1b[0m" }
pub fn on_gray9(input string) string { return "\x1b[48;2;22;22;22m${input}\x1b[0m" }
pub fn on_gray10(input string) string { return "\x1b[48;2;25;25;25m${input}\x1b[0m" }
pub fn on_gray11(input string) string { return "\x1b[48;2;28;28;28m${input}\x1b[0m" }
pub fn on_gray12(input string) string { return "\x1b[48;2;30;30;30m${input}\x1b[0m" }
pub fn on_gray13(input string) string { return "\x1b[48;2;30;30;30m${input}\x1b[0m" }
pub fn on_gray14(input string) string { return "\x1b[48;2;35;35;35m${input}\x1b[0m" }
pub fn on_gray15(input string) string { return "\x1b[48;2;35;35;35m${input}\x1b[0m" }
pub fn on_gray16(input string) string { return "\x1b[48;2;40;40;40m${input}\x1b[0m" }
pub fn on_gray17(input string) string { return "\x1b[48;2;40;40;40m${input}\x1b[0m" }
pub fn on_gray18(input string) string { return "\x1b[48;2;45;45;45m${input}\x1b[0m" }
pub fn on_gray19(input string) string { return "\x1b[48;2;45;45;45m${input}\x1b[0m" }
pub fn on_gray20(input string) string { return "\x1b[48;2;51;51;51m${input}\x1b[0m" }
pub fn on_gray21(input string) string { return "\x1b[48;2;53;53;53m${input}\x1b[0m" }
pub fn on_gray22(input string) string { return "\x1b[48;2;56;56;56m${input}\x1b[0m" }
pub fn on_gray23(input string) string { return "\x1b[48;2;58;58;58m${input}\x1b[0m" }
pub fn on_gray24(input string) string { return "\x1b[48;2;58;58;58m${input}\x1b[0m" }
pub fn on_gray25(input string) string { return "\x1b[48;2;63;63;63m${input}\x1b[0m" }
pub fn on_gray26(input string) string { return "\x1b[48;2;63;63;63m${input}\x1b[0m" }
pub fn on_gray27(input string) string { return "\x1b[48;2;68;68;68m${input}\x1b[0m" }
pub fn on_gray28(input string) string { return "\x1b[48;2;68;68;68m${input}\x1b[0m" }
pub fn on_gray29(input string) string { return "\x1b[48;2;73;73;73m${input}\x1b[0m" }
pub fn on_gray30(input string) string { return "\x1b[48;2;76;76;76m${input}\x1b[0m" }
pub fn on_gray31(input string) string { return "\x1b[48;2;79;79;79m${input}\x1b[0m" }
pub fn on_gray32(input string) string { return "\x1b[48;2;81;81;81m${input}\x1b[0m" }
pub fn on_gray33(input string) string { return "\x1b[48;2;81;81;81m${input}\x1b[0m" }
pub fn on_gray34(input string) string { return "\x1b[48;2;86;86;86m${input}\x1b[0m" }
pub fn on_gray35(input string) string { return "\x1b[48;2;86;86;86m${input}\x1b[0m" }
pub fn on_gray36(input string) string { return "\x1b[48;2;91;91;91m${input}\x1b[0m" }
pub fn on_gray37(input string) string { return "\x1b[48;2;91;91;91m${input}\x1b[0m" }
pub fn on_gray38(input string) string { return "\x1b[48;2;96;96;96m${input}\x1b[0m" }
pub fn on_gray39(input string) string { return "\x1b[48;2;96;96;96m${input}\x1b[0m" }
pub fn on_gray40(input string) string { return "\x1b[48;2;102;102;102m${input}\x1b[0m" }
pub fn on_dimgray(input string) string { return "\x1b[48;2;104;104;104m${input}\x1b[0m" }
pub fn on_gray42(input string) string { return "\x1b[48;2;107;107;107m${input}\x1b[0m" }
pub fn on_gray43(input string) string { return "\x1b[48;2;109;109;109m${input}\x1b[0m" }
pub fn on_gray44(input string) string { return "\x1b[48;2;109;109;109m${input}\x1b[0m" }
pub fn on_gray45(input string) string { return "\x1b[48;2;114;114;114m${input}\x1b[0m" }
pub fn on_gray46(input string) string { return "\x1b[48;2;114;114;114m${input}\x1b[0m" }
pub fn on_gray47(input string) string { return "\x1b[48;2;119;119;119m${input}\x1b[0m" }
pub fn on_gray48(input string) string { return "\x1b[48;2;119;119;119m${input}\x1b[0m" }
pub fn on_gray49(input string) string { return "\x1b[48;2;124;124;124m${input}\x1b[0m" }
pub fn on_gray50(input string) string { return "\x1b[48;2;124;124;124m${input}\x1b[0m" }
pub fn on_webgray(input string) string { return "\x1b[48;2;127;127;127m${input}\x1b[0m" }
pub fn on_gray51(input string) string { return "\x1b[48;2;130;130;130m${input}\x1b[0m" }
pub fn on_gray52(input string) string { return "\x1b[48;2;132;132;132m${input}\x1b[0m" }
pub fn on_gray53(input string) string { return "\x1b[48;2;132;132;132m${input}\x1b[0m" }
pub fn on_gray54(input string) string { return "\x1b[48;2;137;137;137m${input}\x1b[0m" }
pub fn on_gray55(input string) string { return "\x1b[48;2;137;137;137m${input}\x1b[0m" }
pub fn on_gray56(input string) string { return "\x1b[48;2;142;142;142m${input}\x1b[0m" }
pub fn on_gray57(input string) string { return "\x1b[48;2;142;142;142m${input}\x1b[0m" }
pub fn on_gray58(input string) string { return "\x1b[48;2;147;147;147m${input}\x1b[0m" }
pub fn on_gray59(input string) string { return "\x1b[48;2;147;147;147m${input}\x1b[0m" }
pub fn on_gray60(input string) string { return "\x1b[48;2;153;153;153m${input}\x1b[0m" }
pub fn on_gray61(input string) string { return "\x1b[48;2;155;155;155m${input}\x1b[0m" }
pub fn on_gray62(input string) string { return "\x1b[48;2;158;158;158m${input}\x1b[0m" }
pub fn on_gray63(input string) string { return "\x1b[48;2;160;160;160m${input}\x1b[0m" }
pub fn on_gray64(input string) string { return "\x1b[48;2;160;160;160m${input}\x1b[0m" }
pub fn on_gray65(input string) string { return "\x1b[48;2;165;165;165m${input}\x1b[0m" }
pub fn on_gray66(input string) string { return "\x1b[48;2;165;165;165m${input}\x1b[0m" }
pub fn on_darkgray(input string) string { return "\x1b[48;2;168;168;168m${input}\x1b[0m" }
pub fn on_gray67(input string) string { return "\x1b[48;2;170;170;170m${input}\x1b[0m" }
pub fn on_gray68(input string) string { return "\x1b[48;2;170;170;170m${input}\x1b[0m" }
pub fn on_gray69(input string) string { return "\x1b[48;2;175;175;175m${input}\x1b[0m" }
pub fn on_gray70(input string) string { return "\x1b[48;2;178;178;178m${input}\x1b[0m" }
pub fn on_gray71(input string) string { return "\x1b[48;2;181;181;181m${input}\x1b[0m" }
pub fn on_gray72(input string) string { return "\x1b[48;2;183;183;183m${input}\x1b[0m" }
pub fn on_gray73(input string) string { return "\x1b[48;2;183;183;183m${input}\x1b[0m" }
pub fn on_gray74(input string) string { return "\x1b[48;2;188;188;188m${input}\x1b[0m" }
pub fn on_gray(input string) string { return "\x1b[48;2;188;188;188m${input}\x1b[0m" }
pub fn on_gray75(input string) string { return "\x1b[48;2;188;188;188m${input}\x1b[0m" }
pub fn on_silver(input string) string { return "\x1b[48;2;191;191;191m${input}\x1b[0m" }
pub fn on_gray76(input string) string { return "\x1b[48;2;193;193;193m${input}\x1b[0m" }
pub fn on_gray77(input string) string { return "\x1b[48;2;193;193;193m${input}\x1b[0m" }
pub fn on_gray78(input string) string { return "\x1b[48;2;198;198;198m${input}\x1b[0m" }
pub fn on_gray79(input string) string { return "\x1b[48;2;198;198;198m${input}\x1b[0m" }
pub fn on_gray80(input string) string { return "\x1b[48;2;204;204;204m${input}\x1b[0m" }
pub fn on_gray81(input string) string { return "\x1b[48;2;206;206;206m${input}\x1b[0m" }
pub fn on_gray82(input string) string { return "\x1b[48;2;209;209;209m${input}\x1b[0m" }
pub fn on_lightgray(input string) string { return "\x1b[48;2;209;209;209m${input}\x1b[0m" }
pub fn on_gray83(input string) string { return "\x1b[48;2;211;211;211m${input}\x1b[0m" }
pub fn on_gray84(input string) string { return "\x1b[48;2;211;211;211m${input}\x1b[0m" }
pub fn on_gray85(input string) string { return "\x1b[48;2;216;216;216m${input}\x1b[0m" }
pub fn on_gray86(input string) string { return "\x1b[48;2;216;216;216m${input}\x1b[0m" }
pub fn on_gainsboro(input string) string { return "\x1b[48;2;219;219;219m${input}\x1b[0m" }
pub fn on_gray87(input string) string { return "\x1b[48;2;221;221;221m${input}\x1b[0m" }
pub fn on_gray88(input string) string { return "\x1b[48;2;221;221;221m${input}\x1b[0m" }
pub fn on_gray89(input string) string { return "\x1b[48;2;226;226;226m${input}\x1b[0m" }
pub fn on_gray90(input string) string { return "\x1b[48;2;226;226;226m${input}\x1b[0m" }
pub fn on_gray91(input string) string { return "\x1b[48;2;232;232;232m${input}\x1b[0m" }
pub fn on_gray92(input string) string { return "\x1b[48;2;234;234;234m${input}\x1b[0m" }
pub fn on_gray93(input string) string { return "\x1b[48;2;234;234;234m${input}\x1b[0m" }
pub fn on_gray94(input string) string { return "\x1b[48;2;239;239;239m${input}\x1b[0m" }
pub fn on_gray95(input string) string { return "\x1b[48;2;239;239;239m${input}\x1b[0m" }
pub fn on_gray96(input string) string { return "\x1b[48;2;244;244;244m${input}\x1b[0m" }
pub fn on_gray97(input string) string { return "\x1b[48;2;244;244;244m${input}\x1b[0m" }
pub fn on_gray98(input string) string { return "\x1b[48;2;249;249;249m${input}\x1b[0m" }
pub fn on_gray99(input string) string { return "\x1b[48;2;249;249;249m${input}\x1b[0m" }
pub fn on_gray100(input string) string { return "\x1b[48;2;255;255;255m${input}\x1b[0m" }
